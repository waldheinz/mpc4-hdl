
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- This file was generated with hex2rom written by Daniel Wallner

entity U2732 is
	Port ( A 		: in  STD_LOGIC_VECTOR (11 downto 0);
           CE_n 	: in  STD_LOGIC;
           OE_n	: in  STD_LOGIC;
           D 		: out STD_LOGIC_VECTOR (7 downto 0));
end U2732;

architecture rtl of U2732 is
	subtype ROM_WORD is std_logic_vector(7 downto 0);
	type ROM_TABLE is array(0 to 4095) of ROM_WORD;
	constant ROM: ROM_TABLE := ROM_TABLE'(
		"11110011",	-- 0x0000
		"11000011",	-- 0x0001
		"00010011",	-- 0x0002
		"11000000",	-- 0x0003
		"11000011",	-- 0x0004
		"00011010",	-- 0x0005
		"11000100",	-- 0x0006
		"11000011",	-- 0x0007
		"11100110",	-- 0x0008
		"11111100",	-- 0x0009
		"11000011",	-- 0x000A
		"00110100",	-- 0x000B
		"11000100",	-- 0x000C
		"11000011",	-- 0x000D
		"00111110",	-- 0x000E
		"11000100",	-- 0x000F
		"11000011",	-- 0x0010
		"10010101",	-- 0x0011
		"11000000",	-- 0x0012
		"00111110",	-- 0x0013
		"11001111",	-- 0x0014
		"11010011",	-- 0x0015
		"11101110",	-- 0x0016
		"00111110",	-- 0x0017
		"10000000",	-- 0x0018
		"11010011",	-- 0x0019
		"11101110",	-- 0x001A
		"00111110",	-- 0x001B
		"01000000",	-- 0x001C
		"11010011",	-- 0x001D
		"11101100",	-- 0x001E
		"11000011",	-- 0x001F
		"01001111",	-- 0x0020
		"11000000",	-- 0x0021
		"11000011",	-- 0x0022
		"10111001",	-- 0x0023
		"11000101",	-- 0x0024
		"11011011",	-- 0x0025
		"11111110",	-- 0x0026
		"01111110",	-- 0x0027
		"11010011",	-- 0x0028
		"11111110",	-- 0x0029
		"11001001",	-- 0x002A
		"11011011",	-- 0x002B
		"11111110",	-- 0x002C
		"01110001",	-- 0x002D
		"11010011",	-- 0x002E
		"11111110",	-- 0x002F
		"11001001",	-- 0x0030
		"11000011",	-- 0x0031
		"10111110",	-- 0x0032
		"11000011",	-- 0x0033
		"01001111",	-- 0x0034
		"11000011",	-- 0x0035
		"11000101",	-- 0x0036
		"11000101",	-- 0x0037
		"11000011",	-- 0x0038
		"00011101",	-- 0x0039
		"11000100",	-- 0x003A
		"00001101",	-- 0x003B
		"01001101",	-- 0x003C
		"01001111",	-- 0x003D
		"01001110",	-- 0x003E
		"01001001",	-- 0x003F
		"00100000",	-- 0x0040
		"01001101",	-- 0x0041
		"01010000",	-- 0x0042
		"01000011",	-- 0x0043
		"00100000",	-- 0x0044
		"01010110",	-- 0x0045
		"00101110",	-- 0x0046
		"00110000",	-- 0x0047
		"00110001",	-- 0x0048
		"00001101",	-- 0x0049
		"00001101",	-- 0x004A
		"01001001",	-- 0x004B
		"01001110",	-- 0x004C
		"01001001",	-- 0x004D
		"01010100",	-- 0x004E
		"00100001",	-- 0x004F
		"01011010",	-- 0x0050
		"11111100",	-- 0x0051
		"00000110",	-- 0x0052
		"10000010",	-- 0x0053
		"10101111",	-- 0x0054
		"01110111",	-- 0x0055
		"00100011",	-- 0x0056
		"00010000",	-- 0x0057
		"11111011",	-- 0x0058
		"00110001",	-- 0x0059
		"11011100",	-- 0x005A
		"11111100",	-- 0x005B
		"11001101",	-- 0x005C
		"11101111",	-- 0x005D
		"11000011",	-- 0x005E
		"00100001",	-- 0x005F
		"00100010",	-- 0x0060
		"11000000",	-- 0x0061
		"00010001",	-- 0x0062
		"11100110",	-- 0x0063
		"11111100",	-- 0x0064
		"00000001",	-- 0x0065
		"00011001",	-- 0x0066
		"00000000",	-- 0x0067
		"11101101",	-- 0x0068
		"10110000",	-- 0x0069
		"00100001",	-- 0x006A
		"10110000",	-- 0x006B
		"11000101",	-- 0x006C
		"00010001",	-- 0x006D
		"11011100",	-- 0x006E
		"11111100",	-- 0x006F
		"00000001",	-- 0x0070
		"00001001",	-- 0x0071
		"00000000",	-- 0x0072
		"11101101",	-- 0x0073
		"10110000",	-- 0x0074
		"00100001",	-- 0x0075
		"01001010",	-- 0x0076
		"11000000",	-- 0x0077
		"00000110",	-- 0x0078
		"00000101",	-- 0x0079
		"11001101",	-- 0x007A
		"00111100",	-- 0x007B
		"11000011",	-- 0x007C
		"00111110",	-- 0x007D
		"11000011",	-- 0x007E
		"00100001",	-- 0x007F
		"10010101",	-- 0x0080
		"11000000",	-- 0x0081
		"00110010",	-- 0x0082
		"00111000",	-- 0x0083
		"00000000",	-- 0x0084
		"00100010",	-- 0x0085
		"00111001",	-- 0x0086
		"00000000",	-- 0x0087
		"00111110",	-- 0x0088
		"10000001",	-- 0x0089
		"00110010",	-- 0x008A
		"01011011",	-- 0x008B
		"11111100",	-- 0x008C
		"00100001",	-- 0x008D
		"00000000",	-- 0x008E
		"00000000",	-- 0x008F
		"00111110",	-- 0x0090
		"11111101",	-- 0x0091
		"11101101",	-- 0x0092
		"01000111",	-- 0x0093
		"11100101",	-- 0x0094
		"11110011",	-- 0x0095
		"11101101",	-- 0x0096
		"01011110",	-- 0x0097
		"00100010",	-- 0x0098
		"01001110",	-- 0x0099
		"11111100",	-- 0x009A
		"11100001",	-- 0x009B
		"00100010",	-- 0x009C
		"01010110",	-- 0x009D
		"11111100",	-- 0x009E
		"11101101",	-- 0x009F
		"01110011",	-- 0x00A0
		"01011000",	-- 0x00A1
		"11111100",	-- 0x00A2
		"00110001",	-- 0x00A3
		"01010110",	-- 0x00A4
		"11111100",	-- 0x00A5
		"11110101",	-- 0x00A6
		"11000101",	-- 0x00A7
		"11010101",	-- 0x00A8
		"00001000",	-- 0x00A9
		"11011001",	-- 0x00AA
		"00111011",	-- 0x00AB
		"00111011",	-- 0x00AC
		"11110101",	-- 0x00AD
		"11000101",	-- 0x00AE
		"11010101",	-- 0x00AF
		"11100101",	-- 0x00B0
		"11011101",	-- 0x00B1
		"11100101",	-- 0x00B2
		"11111101",	-- 0x00B3
		"11100101",	-- 0x00B4
		"11101101",	-- 0x00B5
		"01010111",	-- 0x00B6
		"11110101",	-- 0x00B7
		"00111110",	-- 0x00B8
		"11111101",	-- 0x00B9
		"11101101",	-- 0x00BA
		"01000111",	-- 0x00BB
		"00111010",	-- 0x00BC
		"01011011",	-- 0x00BD
		"11111100",	-- 0x00BE
		"11001011",	-- 0x00BF
		"11000111",	-- 0x00C0
		"00110010",	-- 0x00C1
		"01011011",	-- 0x00C2
		"11111100",	-- 0x00C3
		"00110001",	-- 0x00C4
		"10011110",	-- 0x00C5
		"11111100",	-- 0x00C6
		"11111011",	-- 0x00C7
		"00100001",	-- 0x00C8
		"00111011",	-- 0x00C9
		"11000000",	-- 0x00CA
		"00000110",	-- 0x00CB
		"00001111",	-- 0x00CC
		"11001101",	-- 0x00CD
		"00111100",	-- 0x00CE
		"11000011",	-- 0x00CF
		"00100001",	-- 0x00D0
		"01011011",	-- 0x00D1
		"11111100",	-- 0x00D2
		"11001011",	-- 0x00D3
		"01111110",	-- 0x00D4
		"11001011",	-- 0x00D5
		"10111110",	-- 0x00D6
		"11000010",	-- 0x00D7
		"00110110",	-- 0x00D8
		"11000101",	-- 0x00D9
		"00111110",	-- 0x00DA
		"00111010",	-- 0x00DB
		"11001101",	-- 0x00DC
		"00110111",	-- 0x00DD
		"11000001",	-- 0x00DE
		"11001101",	-- 0x00DF
		"00011111",	-- 0x00E0
		"11000001",	-- 0x00E1
		"11001101",	-- 0x00E2
		"11100000",	-- 0x00E3
		"11000011",	-- 0x00E4
		"00100001",	-- 0x00E5
		"00000100",	-- 0x00E6
		"11000001",	-- 0x00E7
		"00000001",	-- 0x00E8
		"00001001",	-- 0x00E9
		"00000000",	-- 0x00EA
		"11101101",	-- 0x00EB
		"10110001",	-- 0x00EC
		"00100000",	-- 0x00ED
		"00001010",	-- 0x00EE
		"00100001",	-- 0x00EF
		"00001101",	-- 0x00F0
		"11000001",	-- 0x00F1
		"00001001",	-- 0x00F2
		"00001001",	-- 0x00F3
		"01111110",	-- 0x00F4
		"00100011",	-- 0x00F5
		"01100110",	-- 0x00F6
		"01101111",	-- 0x00F7
		"11101001",	-- 0x00F8
		"00110001",	-- 0x00F9
		"10011110",	-- 0x00FA
		"11111100",	-- 0x00FB
		"00111110",	-- 0x00FC
		"00111111",	-- 0x00FD
		"11001101",	-- 0x00FE
		"00110111",	-- 0x00FF
		"11000001",	-- 0x0100
		"11000011",	-- 0x0101
		"01100001",	-- 0x0102
		"11000010",	-- 0x0103
		"01001100",	-- 0x0104
		"01001001",	-- 0x0105
		"01001111",	-- 0x0106
		"01000111",	-- 0x0107
		"01000100",	-- 0x0108
		"01000110",	-- 0x0109
		"01001101",	-- 0x010A
		"01010011",	-- 0x010B
		"01011000",	-- 0x010C
		"11001110",	-- 0x010D
		"11000010",	-- 0x010E
		"10100000",	-- 0x010F
		"11000010",	-- 0x0110
		"10000110",	-- 0x0111
		"11000010",	-- 0x0112
		"01110111",	-- 0x0113
		"11000010",	-- 0x0114
		"00001011",	-- 0x0115
		"11000010",	-- 0x0116
		"10001101",	-- 0x0117
		"11000011",	-- 0x0118
		"11010111",	-- 0x0119
		"11000011",	-- 0x011A
		"11001100",	-- 0x011B
		"11000011",	-- 0x011C
		"00110110",	-- 0x011D
		"11000101",	-- 0x011E
		"11000101",	-- 0x011F
		"11010101",	-- 0x0120
		"11001101",	-- 0x0121
		"01001110",	-- 0x0122
		"11000001",	-- 0x0123
		"11001101",	-- 0x0124
		"01000001",	-- 0x0125
		"11000001",	-- 0x0126
		"11010001",	-- 0x0127
		"11000001",	-- 0x0128
		"11001001",	-- 0x0129
		"00011010",	-- 0x012A
		"11110101",	-- 0x012B
		"00001111",	-- 0x012C
		"00001111",	-- 0x012D
		"00001111",	-- 0x012E
		"00001111",	-- 0x012F
		"11001101",	-- 0x0130
		"00110100",	-- 0x0131
		"11000001",	-- 0x0132
		"11110001",	-- 0x0133
		"11001101",	-- 0x0134
		"01010111",	-- 0x0135
		"11000001",	-- 0x0136
		"11110101",	-- 0x0137
		"11000101",	-- 0x0138
		"11010101",	-- 0x0139
		"11001101",	-- 0x013A
		"01000001",	-- 0x013B
		"11000001",	-- 0x013C
		"11010001",	-- 0x013D
		"11000001",	-- 0x013E
		"11110001",	-- 0x013F
		"11001001",	-- 0x0140
		"11001101",	-- 0x0141
		"00110100",	-- 0x0142
		"11000100",	-- 0x0143
		"11111110",	-- 0x0144
		"00001101",	-- 0x0145
		"11110101",	-- 0x0146
		"00111110",	-- 0x0147
		"00001010",	-- 0x0148
		"11001100",	-- 0x0149
		"00110100",	-- 0x014A
		"11000100",	-- 0x014B
		"11110001",	-- 0x014C
		"11001001",	-- 0x014D
		"11001101",	-- 0x014E
		"00011010",	-- 0x014F
		"11000100",	-- 0x0150
		"11111110",	-- 0x0151
		"00001101",	-- 0x0152
		"11000000",	-- 0x0153
		"11110101",	-- 0x0154
		"00011000",	-- 0x0155
		"11110010",	-- 0x0156
		"11100110",	-- 0x0157
		"00001111",	-- 0x0158
		"11000110",	-- 0x0159
		"00110000",	-- 0x015A
		"11111110",	-- 0x015B
		"00111010",	-- 0x015C
		"11111000",	-- 0x015D
		"11000110",	-- 0x015E
		"00000111",	-- 0x015F
		"11001001",	-- 0x0160
		"11010110",	-- 0x0161
		"00110000",	-- 0x0162
		"11111110",	-- 0x0163
		"00001010",	-- 0x0164
		"11111000",	-- 0x0165
		"11010110",	-- 0x0166
		"00000111",	-- 0x0167
		"11001001",	-- 0x0168
		"01111001",	-- 0x0169
		"11111110",	-- 0x016A
		"00110000",	-- 0x016B
		"00111111",	-- 0x016C
		"11010000",	-- 0x016D
		"11111110",	-- 0x016E
		"00111010",	-- 0x016F
		"11011000",	-- 0x0170
		"11111110",	-- 0x0171
		"01000001",	-- 0x0172
		"00111111",	-- 0x0173
		"11010000",	-- 0x0174
		"11111110",	-- 0x0175
		"01000111",	-- 0x0176
		"11001001",	-- 0x0177
		"11111110",	-- 0x0178
		"00110000",	-- 0x0179
		"00111111",	-- 0x017A
		"11010000",	-- 0x017B
		"11111110",	-- 0x017C
		"00111010",	-- 0x017D
		"11001001",	-- 0x017E
		"01111001",	-- 0x017F
		"11111110",	-- 0x0180
		"00101100",	-- 0x0181
		"00110111",	-- 0x0182
		"11001000",	-- 0x0183
		"11111110",	-- 0x0184
		"00100000",	-- 0x0185
		"00110111",	-- 0x0186
		"11001000",	-- 0x0187
		"11111110",	-- 0x0188
		"00001101",	-- 0x0189
		"00110111",	-- 0x018A
		"11001000",	-- 0x018B
		"00111111",	-- 0x018C
		"11001001",	-- 0x018D
		"11100101",	-- 0x018E
		"10110111",	-- 0x018F
		"11101101",	-- 0x0190
		"01010010",	-- 0x0191
		"00111111",	-- 0x0192
		"11100001",	-- 0x0193
		"11001001",	-- 0x0194
		"11100101",	-- 0x0195
		"00100001",	-- 0x0196
		"00000000",	-- 0x0197
		"00000000",	-- 0x0198
		"01011100",	-- 0x0199
		"11001101",	-- 0x019A
		"00011111",	-- 0x019B
		"11000001",	-- 0x019C
		"11001101",	-- 0x019D
		"11100000",	-- 0x019E
		"11000011",	-- 0x019F
		"01001111",	-- 0x01A0
		"11001101",	-- 0x01A1
		"01111111",	-- 0x01A2
		"11000001",	-- 0x01A3
		"00110000",	-- 0x01A4
		"00001001",	-- 0x01A5
		"01010001",	-- 0x01A6
		"11100101",	-- 0x01A7
		"11000001",	-- 0x01A8
		"11100001",	-- 0x01A9
		"01111011",	-- 0x01AA
		"10110111",	-- 0x01AB
		"11001000",	-- 0x01AC
		"00110111",	-- 0x01AD
		"11001001",	-- 0x01AE
		"11001101",	-- 0x01AF
		"01101001",	-- 0x01B0
		"11000001",	-- 0x01B1
		"11010010",	-- 0x01B2
		"11111001",	-- 0x01B3
		"11000000",	-- 0x01B4
		"01111001",	-- 0x01B5
		"11001101",	-- 0x01B6
		"01100001",	-- 0x01B7
		"11000001",	-- 0x01B8
		"00011110",	-- 0x01B9
		"11111111",	-- 0x01BA
		"00101001",	-- 0x01BB
		"00101001",	-- 0x01BC
		"00101001",	-- 0x01BD
		"00101001",	-- 0x01BE
		"00000110",	-- 0x01BF
		"00000000",	-- 0x01C0
		"01001111",	-- 0x01C1
		"00001001",	-- 0x01C2
		"00011000",	-- 0x01C3
		"11010101",	-- 0x01C4
		"01111100",	-- 0x01C5
		"11001101",	-- 0x01C6
		"00101011",	-- 0x01C7
		"11000001",	-- 0x01C8
		"01111101",	-- 0x01C9
		"11000011",	-- 0x01CA
		"00101011",	-- 0x01CB
		"11000001",	-- 0x01CC
		"00101110",	-- 0x01CD
		"00000011",	-- 0x01CE
		"01111001",	-- 0x01CF
		"11100110",	-- 0x01D0
		"00000011",	-- 0x01D1
		"01100111",	-- 0x01D2
		"11001101",	-- 0x01D3
		"10010101",	-- 0x01D4
		"11000001",	-- 0x01D5
		"11010010",	-- 0x01D6
		"11111001",	-- 0x01D7
		"11000000",	-- 0x01D8
		"11000101",	-- 0x01D9
		"00101101",	-- 0x01DA
		"00100101",	-- 0x01DB
		"01111010",	-- 0x01DC
		"00101000",	-- 0x01DD
		"00001010",	-- 0x01DE
		"11111110",	-- 0x01DF
		"00001101",	-- 0x01E0
		"11001010",	-- 0x01E1
		"11111001",	-- 0x01E2
		"11000000",	-- 0x01E3
		"00110010",	-- 0x01E4
		"01011100",	-- 0x01E5
		"11111100",	-- 0x01E6
		"00011000",	-- 0x01E7
		"11101010",	-- 0x01E8
		"11111110",	-- 0x01E9
		"00001101",	-- 0x01EA
		"11000010",	-- 0x01EB
		"11111001",	-- 0x01EC
		"11000000",	-- 0x01ED
		"00000001",	-- 0x01EE
		"11111111",	-- 0x01EF
		"11111111",	-- 0x01F0
		"01111101",	-- 0x01F1
		"10110111",	-- 0x01F2
		"00101000",	-- 0x01F3
		"00000100",	-- 0x01F4
		"11000101",	-- 0x01F5
		"00101101",	-- 0x01F6
		"00100000",	-- 0x01F7
		"11111100",	-- 0x01F8
		"11000001",	-- 0x01F9
		"11010001",	-- 0x01FA
		"11100001",	-- 0x01FB
		"11001101",	-- 0x01FC
		"10001110",	-- 0x01FD
		"11000001",	-- 0x01FE
		"00110000",	-- 0x01FF
		"00000000",	-- 0x0200
		"11100011",	-- 0x0201
		"11010101",	-- 0x0202
		"11000101",	-- 0x0203
		"11100101",	-- 0x0204
		"00111101",	-- 0x0205
		"11111000",	-- 0x0206
		"11100001",	-- 0x0207
		"11100011",	-- 0x0208
		"00011000",	-- 0x0209
		"11111010",	-- 0x020A
		"11001101",	-- 0x020B
		"01100111",	-- 0x020C
		"11000010",	-- 0x020D
		"11000101",	-- 0x020E
		"11000001",	-- 0x020F
		"00000110",	-- 0x0210
		"00000000",	-- 0x0211
		"11100101",	-- 0x0212
		"11001101",	-- 0x0213
		"11000101",	-- 0x0214
		"11000001",	-- 0x0215
		"10101111",	-- 0x0216
		"10110000",	-- 0x0217
		"11000100",	-- 0x0218
		"01000100",	-- 0x0219
		"11000011",	-- 0x021A
		"11001101",	-- 0x021B
		"01000100",	-- 0x021C
		"11000011",	-- 0x021D
		"11001101",	-- 0x021E
		"11101001",	-- 0x021F
		"11111100",	-- 0x0220
		"00100000",	-- 0x0221
		"00100000",	-- 0x0222
		"11001101",	-- 0x0223
		"00101011",	-- 0x0224
		"11000001",	-- 0x0225
		"11001101",	-- 0x0226
		"10001110",	-- 0x0227
		"11000001",	-- 0x0228
		"00111000",	-- 0x0229
		"00101010",	-- 0x022A
		"00100011",	-- 0x022B
		"01111101",	-- 0x022C
		"11100110",	-- 0x022D
		"00001111",	-- 0x022E
		"00100000",	-- 0x022F
		"11100101",	-- 0x0230
		"11001101",	-- 0x0231
		"01001000",	-- 0x0232
		"11000011",	-- 0x0233
		"00111010",	-- 0x0234
		"01011100",	-- 0x0235
		"11111100",	-- 0x0236
		"11111110",	-- 0x0237
		"00101100",	-- 0x0238
		"00100000",	-- 0x0239
		"11011000",	-- 0x023A
		"10101111",	-- 0x023B
		"10110000",	-- 0x023C
		"00100000",	-- 0x023D
		"11010000",	-- 0x023E
		"00000100",	-- 0x023F
		"11100001",	-- 0x0240
		"00011000",	-- 0x0241
		"11001111",	-- 0x0242
		"11111110",	-- 0x0243
		"00100000",	-- 0x0244
		"00111000",	-- 0x0245
		"00001001",	-- 0x0246
		"11111110",	-- 0x0247
		"01111111",	-- 0x0248
		"00110000",	-- 0x0249
		"00000101",	-- 0x024A
		"11001101",	-- 0x024B
		"00110111",	-- 0x024C
		"11000001",	-- 0x024D
		"00011000",	-- 0x024E
		"11010110",	-- 0x024F
		"11001101",	-- 0x0250
		"01000100",	-- 0x0251
		"11000011",	-- 0x0252
		"00011000",	-- 0x0253
		"11010001",	-- 0x0254
		"00111010",	-- 0x0255
		"01011100",	-- 0x0256
		"11111100",	-- 0x0257
		"11111110",	-- 0x0258
		"00101100",	-- 0x0259
		"00100000",	-- 0x025A
		"00000100",	-- 0x025B
		"10101111",	-- 0x025C
		"10110000",	-- 0x025D
		"00101000",	-- 0x025E
		"11010001",	-- 0x025F
		"11100001",	-- 0x0260
		"11001101",	-- 0x0261
		"01001000",	-- 0x0262
		"11000011",	-- 0x0263
		"11000011",	-- 0x0264
		"11011010",	-- 0x0265
		"11000000",	-- 0x0266
		"00001110",	-- 0x0267
		"00000010",	-- 0x0268
		"11001101",	-- 0x0269
		"11001101",	-- 0x026A
		"11000001",	-- 0x026B
		"11010001",	-- 0x026C
		"11100001",	-- 0x026D
		"11001001",	-- 0x026E
		"00001110",	-- 0x026F
		"00000011",	-- 0x0270
		"11001101",	-- 0x0271
		"11001101",	-- 0x0272
		"11000001",	-- 0x0273
		"11000001",	-- 0x0274
		"00011000",	-- 0x0275
		"11110101",	-- 0x0276
		"11001101",	-- 0x0277
		"01101111",	-- 0x0278
		"11000010",	-- 0x0279
		"11001101",	-- 0x027A
		"11101111",	-- 0x027B
		"11111100",	-- 0x027C
		"11001101",	-- 0x027D
		"10001110",	-- 0x027E
		"11000001",	-- 0x027F
		"11011010",	-- 0x0280
		"11011010",	-- 0x0281
		"11000000",	-- 0x0282
		"00100011",	-- 0x0283
		"00011000",	-- 0x0284
		"11110100",	-- 0x0285
		"11001101",	-- 0x0286
		"01101111",	-- 0x0287
		"11000010",	-- 0x0288
		"11001101",	-- 0x0289
		"11101001",	-- 0x028A
		"11111100",	-- 0x028B
		"11100101",	-- 0x028C
		"11000101",	-- 0x028D
		"01100000",	-- 0x028E
		"01101001",	-- 0x028F
		"01001111",	-- 0x0290
		"11001101",	-- 0x0291
		"11101111",	-- 0x0292
		"11111100",	-- 0x0293
		"11000001",	-- 0x0294
		"11100001",	-- 0x0295
		"00000011",	-- 0x0296
		"11001101",	-- 0x0297
		"10001110",	-- 0x0298
		"11000001",	-- 0x0299
		"00100011",	-- 0x029A
		"00100000",	-- 0x029B
		"11101100",	-- 0x029C
		"11000011",	-- 0x029D
		"11011010",	-- 0x029E
		"11000000",	-- 0x029F
		"11001101",	-- 0x02A0
		"10010101",	-- 0x02A1
		"11000001",	-- 0x02A2
		"11000101",	-- 0x02A3
		"11100001",	-- 0x02A4
		"01111010",	-- 0x02A5
		"11111110",	-- 0x02A6
		"00001101",	-- 0x02A7
		"11001010",	-- 0x02A8
		"11011010",	-- 0x02A9
		"11000000",	-- 0x02AA
		"11001101",	-- 0x02AB
		"11101001",	-- 0x02AC
		"11111100",	-- 0x02AD
		"11001101",	-- 0x02AE
		"00101011",	-- 0x02AF
		"11000001",	-- 0x02B0
		"11001101",	-- 0x02B1
		"10111100",	-- 0x02B2
		"11000010",	-- 0x02B3
		"00110000",	-- 0x02B4
		"00000011",	-- 0x02B5
		"11001101",	-- 0x02B6
		"11101111",	-- 0x02B7
		"11111100",	-- 0x02B8
		"00100011",	-- 0x02B9
		"00011000",	-- 0x02BA
		"11101001",	-- 0x02BB
		"00111110",	-- 0x02BC
		"00101101",	-- 0x02BD
		"11001101",	-- 0x02BE
		"00110111",	-- 0x02BF
		"11000001",	-- 0x02C0
		"11000011",	-- 0x02C1
		"10010101",	-- 0x02C2
		"11000001",	-- 0x02C3
		"00000110",	-- 0x02C4
		"00000010",	-- 0x02C5
		"11001101",	-- 0x02C6
		"00111100",	-- 0x02C7
		"11000011",	-- 0x02C8
		"00111110",	-- 0x02C9
		"00111101",	-- 0x02CA
		"11000011",	-- 0x02CB
		"00110111",	-- 0x02CC
		"11000001",	-- 0x02CD
		"11001101",	-- 0x02CE
		"00011111",	-- 0x02CF
		"11000001",	-- 0x02D0
		"11001101",	-- 0x02D1
		"11100000",	-- 0x02D2
		"11000011",	-- 0x02D3
		"11111110",	-- 0x02D4
		"00001101",	-- 0x02D5
		"00100001",	-- 0x02D6
		"01001101",	-- 0x02D7
		"11000011",	-- 0x02D8
		"00010001",	-- 0x02D9
		"01011001",	-- 0x02DA
		"11111100",	-- 0x02DB
		"00100000",	-- 0x02DC
		"00000110",	-- 0x02DD
		"11001101",	-- 0x02DE
		"00011101",	-- 0x02DF
		"11000011",	-- 0x02E0
		"11000011",	-- 0x02E1
		"11011010",	-- 0x02E2
		"11000000",	-- 0x02E3
		"11111110",	-- 0x02E4
		"00100000",	-- 0x02E5
		"00101000",	-- 0x02E6
		"00000011",	-- 0x02E7
		"11000011",	-- 0x02E8
		"11111001",	-- 0x02E9
		"11000000",	-- 0x02EA
		"11001101",	-- 0x02EB
		"11000100",	-- 0x02EC
		"11000010",	-- 0x02ED
		"11001101",	-- 0x02EE
		"00101010",	-- 0x02EF
		"11000001",	-- 0x02F0
		"11001011",	-- 0x02F1
		"01000110",	-- 0x02F2
		"00101000",	-- 0x02F3
		"00000100",	-- 0x02F4
		"00011011",	-- 0x02F5
		"11001101",	-- 0x02F6
		"00101010",	-- 0x02F7
		"11000001",	-- 0x02F8
		"11010101",	-- 0x02F9
		"11001101",	-- 0x02FA
		"10111100",	-- 0x02FB
		"11000010",	-- 0x02FC
		"01111010",	-- 0x02FD
		"00110000",	-- 0x02FE
		"00001111",	-- 0x02FF
		"11010001",	-- 0x0300
		"11110101",	-- 0x0301
		"01111110",	-- 0x0302
		"11101011",	-- 0x0303
		"01110001",	-- 0x0304
		"11001011",	-- 0x0305
		"01000111",	-- 0x0306
		"00101000",	-- 0x0307
		"00000011",	-- 0x0308
		"00100011",	-- 0x0309
		"01110000",	-- 0x030A
		"00101011",	-- 0x030B
		"11110001",	-- 0x030C
		"11101011",	-- 0x030D
		"11010101",	-- 0x030E
		"11010001",	-- 0x030F
		"00011011",	-- 0x0310
		"00100011",	-- 0x0311
		"11111110",	-- 0x0312
		"00001101",	-- 0x0313
		"00101000",	-- 0x0314
		"11001011",	-- 0x0315
		"10101111",	-- 0x0316
		"10110110",	-- 0x0317
		"11001010",	-- 0x0318
		"01100001",	-- 0x0319
		"11000010",	-- 0x031A
		"00011000",	-- 0x031B
		"11001110",	-- 0x031C
		"01111110",	-- 0x031D
		"10110111",	-- 0x031E
		"11001010",	-- 0x031F
		"01001000",	-- 0x0320
		"11000011",	-- 0x0321
		"11001101",	-- 0x0322
		"11000100",	-- 0x0323
		"11000010",	-- 0x0324
		"11001101",	-- 0x0325
		"00101010",	-- 0x0326
		"11000001",	-- 0x0327
		"11001011",	-- 0x0328
		"01000110",	-- 0x0329
		"00101000",	-- 0x032A
		"00000100",	-- 0x032B
		"00011011",	-- 0x032C
		"11001101",	-- 0x032D
		"00101010",	-- 0x032E
		"11000001",	-- 0x032F
		"00011011",	-- 0x0330
		"11001101",	-- 0x0331
		"01000100",	-- 0x0332
		"11000011",	-- 0x0333
		"11001011",	-- 0x0334
		"01111110",	-- 0x0335
		"11000100",	-- 0x0336
		"01001000",	-- 0x0337
		"11000011",	-- 0x0338
		"00100011",	-- 0x0339
		"00011000",	-- 0x033A
		"11100001",	-- 0x033B
		"01111110",	-- 0x033C
		"11001101",	-- 0x033D
		"00110111",	-- 0x033E
		"11000001",	-- 0x033F
		"00100011",	-- 0x0340
		"00010000",	-- 0x0341
		"11111001",	-- 0x0342
		"11001001",	-- 0x0343
		"00111110",	-- 0x0344
		"00100000",	-- 0x0345
		"00011000",	-- 0x0346
		"00000010",	-- 0x0347
		"00111110",	-- 0x0348
		"00001101",	-- 0x0349
		"11000011",	-- 0x034A
		"00110111",	-- 0x034B
		"11000001",	-- 0x034C
		"01010011",	-- 0x034D
		"01010000",	-- 0x034E
		"00000001",	-- 0x034F
		"01010000",	-- 0x0350
		"01000011",	-- 0x0351
		"10000001",	-- 0x0352
		"01000001",	-- 0x0353
		"00110001",	-- 0x0354
		"00000000",	-- 0x0355
		"01000110",	-- 0x0356
		"00110001",	-- 0x0357
		"00000000",	-- 0x0358
		"01000010",	-- 0x0359
		"00110001",	-- 0x035A
		"00000000",	-- 0x035B
		"01000011",	-- 0x035C
		"00110001",	-- 0x035D
		"00000000",	-- 0x035E
		"01000100",	-- 0x035F
		"00110001",	-- 0x0360
		"00000000",	-- 0x0361
		"01000101",	-- 0x0362
		"00110001",	-- 0x0363
		"00000000",	-- 0x0364
		"01001000",	-- 0x0365
		"00110001",	-- 0x0366
		"00000000",	-- 0x0367
		"01001100",	-- 0x0368
		"00110001",	-- 0x0369
		"10000000",	-- 0x036A
		"01000001",	-- 0x036B
		"00110010",	-- 0x036C
		"00000000",	-- 0x036D
		"01000110",	-- 0x036E
		"00110010",	-- 0x036F
		"00000000",	-- 0x0370
		"01000010",	-- 0x0371
		"00110010",	-- 0x0372
		"00000000",	-- 0x0373
		"01000011",	-- 0x0374
		"00110010",	-- 0x0375
		"00000000",	-- 0x0376
		"01000100",	-- 0x0377
		"00110010",	-- 0x0378
		"00000000",	-- 0x0379
		"01000101",	-- 0x037A
		"00110010",	-- 0x037B
		"00000000",	-- 0x037C
		"01001000",	-- 0x037D
		"00110010",	-- 0x037E
		"00000000",	-- 0x037F
		"01001100",	-- 0x0380
		"00110010",	-- 0x0381
		"10000000",	-- 0x0382
		"01001001",	-- 0x0383
		"01011000",	-- 0x0384
		"00000001",	-- 0x0385
		"01001001",	-- 0x0386
		"01011001",	-- 0x0387
		"00000001",	-- 0x0388
		"01001001",	-- 0x0389
		"01010010",	-- 0x038A
		"00000000",	-- 0x038B
		"00000000",	-- 0x038C
		"11001101",	-- 0x038D
		"10010101",	-- 0x038E
		"11000001",	-- 0x038F
		"11110101",	-- 0x0390
		"01111010",	-- 0x0391
		"11111110",	-- 0x0392
		"00001101",	-- 0x0393
		"11000010",	-- 0x0394
		"11111001",	-- 0x0395
		"11000000",	-- 0x0396
		"11110001",	-- 0x0397
		"00110000",	-- 0x0398
		"00000100",	-- 0x0399
		"11101101",	-- 0x039A
		"01000011",	-- 0x039B
		"01010110",	-- 0x039C
		"11111100",	-- 0x039D
		"11110011",	-- 0x039E
		"00110001",	-- 0x039F
		"01000000",	-- 0x03A0
		"11111100",	-- 0x03A1
		"00111010",	-- 0x03A2
		"01011011",	-- 0x03A3
		"11111100",	-- 0x03A4
		"11001011",	-- 0x03A5
		"10000111",	-- 0x03A6
		"00110010",	-- 0x03A7
		"01011011",	-- 0x03A8
		"11111100",	-- 0x03A9
		"10101111",	-- 0x03AA
		"11110001",	-- 0x03AB
		"11101101",	-- 0x03AC
		"01000111",	-- 0x03AD
		"11111101",	-- 0x03AE
		"11100001",	-- 0x03AF
		"11011101",	-- 0x03B0
		"11100001",	-- 0x03B1
		"11100001",	-- 0x03B2
		"11010001",	-- 0x03B3
		"11000001",	-- 0x03B4
		"11110001",	-- 0x03B5
		"11011001",	-- 0x03B6
		"00001000",	-- 0x03B7
		"11100001",	-- 0x03B8
		"11010001",	-- 0x03B9
		"11000001",	-- 0x03BA
		"11000011",	-- 0x03BB
		"11110101",	-- 0x03BC
		"11111100",	-- 0x03BD
		"11110001",	-- 0x03BE
		"11101101",	-- 0x03BF
		"01111011",	-- 0x03C0
		"01011000",	-- 0x03C1
		"11111100",	-- 0x03C2
		"00101010",	-- 0x03C3
		"01010110",	-- 0x03C4
		"11111100",	-- 0x03C5
		"11100101",	-- 0x03C6
		"00101010",	-- 0x03C7
		"01001110",	-- 0x03C8
		"11111100",	-- 0x03C9
		"11111011",	-- 0x03CA
		"11001001",	-- 0x03CB
		"11001101",	-- 0x03CC
		"10010101",	-- 0x03CD
		"11000001",	-- 0x03CE
		"11101101",	-- 0x03CF
		"01111000",	-- 0x03D0
		"11001101",	-- 0x03D1
		"00101011",	-- 0x03D2
		"11000001",	-- 0x03D3
		"11000011",	-- 0x03D4
		"01100001",	-- 0x03D5
		"11000010",	-- 0x03D6
		"11001101",	-- 0x03D7
		"01100111",	-- 0x03D8
		"11000010",	-- 0x03D9
		"01001101",	-- 0x03DA
		"11101101",	-- 0x03DB
		"01011001",	-- 0x03DC
		"11000011",	-- 0x03DD
		"01100001",	-- 0x03DE
		"11000010",	-- 0x03DF
		"11111110",	-- 0x03E0
		"01000001",	-- 0x03E1
		"11011000",	-- 0x03E2
		"11111110",	-- 0x03E3
		"01011011",	-- 0x03E4
		"11011000",	-- 0x03E5
		"11111110",	-- 0x03E6
		"01100001",	-- 0x03E7
		"11011000",	-- 0x03E8
		"11111110",	-- 0x03E9
		"01111011",	-- 0x03EA
		"11010000",	-- 0x03EB
		"11001011",	-- 0x03EC
		"10101111",	-- 0x03ED
		"11001001",	-- 0x03EE
		"00100001",	-- 0x03EF
		"00101010",	-- 0x03F0
		"11000100",	-- 0x03F1
		"00100010",	-- 0x03F2
		"00000000",	-- 0x03F3
		"11111101",	-- 0x03F4
		"11001101",	-- 0x03F5
		"11010001",	-- 0x03F6
		"11000101",	-- 0x03F7
		"10101111",	-- 0x03F8
		"00110010",	-- 0x03F9
		"01011101",	-- 0x03FA
		"11111100",	-- 0x03FB
		"00100001",	-- 0x03FC
		"00001100",	-- 0x03FD
		"11000100",	-- 0x03FE
		"00001110",	-- 0x03FF
		"11100111",	-- 0x0400
		"00000110",	-- 0x0401
		"00001100",	-- 0x0402
		"11101101",	-- 0x0403
		"10110011",	-- 0x0404
		"00000110",	-- 0x0405
		"00000010",	-- 0x0406
		"00001110",	-- 0x0407
		"11110100",	-- 0x0408
		"11101101",	-- 0x0409
		"10110011",	-- 0x040A
		"11001001",	-- 0x040B
		"00000000",	-- 0x040C
		"00011000",	-- 0x040D
		"00000001",	-- 0x040E
		"00011000",	-- 0x040F
		"00000010",	-- 0x0410
		"00000000",	-- 0x0411
		"00000011",	-- 0x0412
		"11000001",	-- 0x0413
		"00000100",	-- 0x0414
		"01000100",	-- 0x0415
		"00000101",	-- 0x0416
		"01101000",	-- 0x0417
		"01000111",	-- 0x0418
		"00001101",	-- 0x0419
		"11000011",	-- 0x041A
		"11111100",	-- 0x041B
		"11111100",	-- 0x041C
		"00111010",	-- 0x041D
		"01011010",	-- 0x041E
		"11111100",	-- 0x041F
		"10110111",	-- 0x0420
		"00101000",	-- 0x0421
		"11110111",	-- 0x0422
		"11110101",	-- 0x0423
		"10101111",	-- 0x0424
		"00110010",	-- 0x0425
		"01011010",	-- 0x0426
		"11111100",	-- 0x0427
		"11110001",	-- 0x0428
		"11001001",	-- 0x0429
		"11110101",	-- 0x042A
		"11011011",	-- 0x042B
		"11100101",	-- 0x042C
		"00110010",	-- 0x042D
		"01011010",	-- 0x042E
		"11111100",	-- 0x042F
		"11110001",	-- 0x0430
		"11111011",	-- 0x0431
		"11101101",	-- 0x0432
		"01001101",	-- 0x0433
		"01001111",	-- 0x0434
		"11110101",	-- 0x0435
		"00111010",	-- 0x0436
		"01011011",	-- 0x0437
		"11111100",	-- 0x0438
		"11001011",	-- 0x0439
		"01001111",	-- 0x043A
		"00100000",	-- 0x043B
		"11111001",	-- 0x043C
		"11110001",	-- 0x043D
		"11000011",	-- 0x043E
		"11111001",	-- 0x043F
		"11111100",	-- 0x0440
		"00100001",	-- 0x0441
		"01011110",	-- 0x0442
		"11111100",	-- 0x0443
		"00010110",	-- 0x0444
		"00000000",	-- 0x0445
		"01000110",	-- 0x0446
		"00100011",	-- 0x0447
		"00001110",	-- 0x0448
		"11111001",	-- 0x0449
		"11001101",	-- 0x044A
		"01101010",	-- 0x044B
		"11000100",	-- 0x044C
		"00100000",	-- 0x044D
		"00010100",	-- 0x044E
		"11101101",	-- 0x044F
		"10100011",	-- 0x0450
		"00100000",	-- 0x0451
		"11110111",	-- 0x0452
		"00100001",	-- 0x0453
		"01101001",	-- 0x0454
		"11111100",	-- 0x0455
		"11001101",	-- 0x0456
		"01101010",	-- 0x0457
		"11000100",	-- 0x0458
		"01111010",	-- 0x0459
		"00110010",	-- 0x045A
		"01101000",	-- 0x045B
		"11111100",	-- 0x045C
		"11001000",	-- 0x045D
		"00010100",	-- 0x045E
		"11101101",	-- 0x045F
		"10100010",	-- 0x0460
		"00011000",	-- 0x0461
		"11110011",	-- 0x0462
		"10101111",	-- 0x0463
		"01010111",	-- 0x0464
		"11001101",	-- 0x0465
		"01010011",	-- 0x0466
		"11000100",	-- 0x0467
		"00110111",	-- 0x0468
		"11001001",	-- 0x0469
		"11011011",	-- 0x046A
		"11111000",	-- 0x046B
		"11001011",	-- 0x046C
		"01111111",	-- 0x046D
		"00101000",	-- 0x046E
		"11111010",	-- 0x046F
		"10100111",	-- 0x0470
		"11001011",	-- 0x0471
		"01110111",	-- 0x0472
		"11001001",	-- 0x0473
		"00100001",	-- 0x0474
		"11011100",	-- 0x0475
		"11111100",	-- 0x0476
		"00100010",	-- 0x0477
		"00100000",	-- 0x0478
		"11111101",	-- 0x0479
		"11011011",	-- 0x047A
		"11101100",	-- 0x047B
		"11110110",	-- 0x047C
		"00000001",	-- 0x047D
		"11010011",	-- 0x047E
		"11101100",	-- 0x047F
		"00000001",	-- 0x0480
		"00000000",	-- 0x0481
		"00010000",	-- 0x0482
		"11000101",	-- 0x0483
		"00100001",	-- 0x0484
		"11001000",	-- 0x0485
		"11000100",	-- 0x0486
		"00010001",	-- 0x0487
		"01011110",	-- 0x0488
		"11111100",	-- 0x0489
		"00000001",	-- 0x048A
		"00000011",	-- 0x048B
		"00000000",	-- 0x048C
		"11101101",	-- 0x048D
		"10110000",	-- 0x048E
		"11001101",	-- 0x048F
		"01000001",	-- 0x0490
		"11000100",	-- 0x0491
		"00111010",	-- 0x0492
		"01101001",	-- 0x0493
		"11111100",	-- 0x0494
		"11000001",	-- 0x0495
		"11001011",	-- 0x0496
		"01101111",	-- 0x0497
		"11000010",	-- 0x0498
		"10100011",	-- 0x0499
		"11000100",	-- 0x049A
		"00001011",	-- 0x049B
		"01111000",	-- 0x049C
		"10110001",	-- 0x049D
		"11001010",	-- 0x049E
		"10100011",	-- 0x049F
		"11000101",	-- 0x04A0
		"00011000",	-- 0x04A1
		"11100000",	-- 0x04A2
		"00100001",	-- 0x04A3
		"11001011",	-- 0x04A4
		"11000100",	-- 0x04A5
		"00010001",	-- 0x04A6
		"01011110",	-- 0x04A7
		"11111100",	-- 0x04A8
		"00000001",	-- 0x04A9
		"00000100",	-- 0x04AA
		"00000000",	-- 0x04AB
		"11101101",	-- 0x04AC
		"10110000",	-- 0x04AD
		"11001101",	-- 0x04AE
		"01000001",	-- 0x04AF
		"11000100",	-- 0x04B0
		"00100001",	-- 0x04B1
		"11001111",	-- 0x04B2
		"11000100",	-- 0x04B3
		"00010001",	-- 0x04B4
		"01011110",	-- 0x04B5
		"11111100",	-- 0x04B6
		"00000001",	-- 0x04B7
		"00000011",	-- 0x04B8
		"00000000",	-- 0x04B9
		"11101101",	-- 0x04BA
		"10110000",	-- 0x04BB
		"11001101",	-- 0x04BC
		"00001010",	-- 0x04BD
		"11000101",	-- 0x04BE
		"00000110",	-- 0x04BF
		"00000110",	-- 0x04C0
		"00111110",	-- 0x04C1
		"11000011",	-- 0x04C2
		"11010011",	-- 0x04C3
		"11111111",	-- 0x04C4
		"00010000",	-- 0x04C5
		"11111100",	-- 0x04C6
		"11001001",	-- 0x04C7
		"00000010",	-- 0x04C8
		"00000100",	-- 0x04C9
		"00000000",	-- 0x04CA
		"00000011",	-- 0x04CB
		"00000011",	-- 0x04CC
		"11110011",	-- 0x04CD
		"11111110",	-- 0x04CE
		"00000010",	-- 0x04CF
		"00000111",	-- 0x04D0
		"00000000",	-- 0x04D1
		"01111001",	-- 0x04D2
		"10000000",	-- 0x04D3
		"10011111",	-- 0x04D4
		"11111111",	-- 0x04D5
		"00010011",	-- 0x04D6
		"01010100",	-- 0x04D7
		"01111100",	-- 0x04D8
		"01101000",	-- 0x04D9
		"10111100",	-- 0x04DA
		"11010101",	-- 0x04DB
		"11111101",	-- 0x04DC
		"00010010",	-- 0x04DD
		"00100000",	-- 0x04DE
		"10001010",	-- 0x04DF
		"11001111",	-- 0x04E0
		"11100000",	-- 0x04E1
		"00001001",	-- 0x04E2
		"01000110",	-- 0x04E3
		"00000000",	-- 0x04E4
		"00000000",	-- 0x04E5
		"00000000",	-- 0x04E6
		"00000001",	-- 0x04E7
		"00000011",	-- 0x04E8
		"00000101",	-- 0x04E9
		"00100101",	-- 0x04EA
		"11111111",	-- 0x04EB
		"00000011",	-- 0x04EC
		"00001111",	-- 0x04ED
		"00000000",	-- 0x04EE
		"00000001",	-- 0x04EF
		"01111001",	-- 0x04F0
		"10000000",	-- 0x04F1
		"10110011",	-- 0x04F2
		"01111111",	-- 0x04F3
		"00001100",	-- 0x04F4
		"01010100",	-- 0x04F5
		"01111100",	-- 0x04F6
		"01101000",	-- 0x04F7
		"10111100",	-- 0x04F8
		"11010101",	-- 0x04F9
		"11111101",	-- 0x04FA
		"00010010",	-- 0x04FB
		"00100000",	-- 0x04FC
		"10001010",	-- 0x04FD
		"11001111",	-- 0x04FE
		"11100000",	-- 0x04FF
		"00001001",	-- 0x0500
		"01000110",	-- 0x0501
		"00000000",	-- 0x0502
		"00000001",	-- 0x0503
		"00000000",	-- 0x0504
		"00000001",	-- 0x0505
		"00000011",	-- 0x0506
		"00000101",	-- 0x0507
		"00100101",	-- 0x0508
		"11111111",	-- 0x0509
		"11001101",	-- 0x050A
		"01000001",	-- 0x050B
		"11000100",	-- 0x050C
		"11011010",	-- 0x050D
		"10100011",	-- 0x050E
		"11000101",	-- 0x050F
		"00111010",	-- 0x0510
		"01101000",	-- 0x0511
		"11111100",	-- 0x0512
		"10110111",	-- 0x0513
		"11000010",	-- 0x0514
		"10100011",	-- 0x0515
		"11000101",	-- 0x0516
		"00111100",	-- 0x0517
		"00110010",	-- 0x0518
		"01011110",	-- 0x0519
		"11111100",	-- 0x051A
		"00111110",	-- 0x051B
		"00001000",	-- 0x051C
		"00110010",	-- 0x051D
		"01011111",	-- 0x051E
		"11111100",	-- 0x051F
		"11001101",	-- 0x0520
		"01000001",	-- 0x0521
		"11000100",	-- 0x0522
		"11011010",	-- 0x0523
		"10100011",	-- 0x0524
		"11000101",	-- 0x0525
		"00111010",	-- 0x0526
		"01101001",	-- 0x0527
		"11111100",	-- 0x0528
		"11111110",	-- 0x0529
		"10000000",	-- 0x052A
		"00101000",	-- 0x052B
		"11110011",	-- 0x052C
		"11100110",	-- 0x052D
		"11100000",	-- 0x052E
		"11111110",	-- 0x052F
		"00100000",	-- 0x0530
		"00001111",	-- 0x0531
		"11001000",	-- 0x0532
		"11000011",	-- 0x0533
		"10100011",	-- 0x0534
		"11000101",	-- 0x0535
		"00000110",	-- 0x0536
		"00001010",	-- 0x0537
		"11000101",	-- 0x0538
		"11001101",	-- 0x0539
		"01110100",	-- 0x053A
		"11000100",	-- 0x053B
		"00100001",	-- 0x053C
		"11010010",	-- 0x053D
		"11000100",	-- 0x053E
		"00001110",	-- 0x053F
		"11111111",	-- 0x0540
		"00000110",	-- 0x0541
		"00010000",	-- 0x0542
		"11101101",	-- 0x0543
		"10110011",	-- 0x0544
		"00100001",	-- 0x0545
		"11100010",	-- 0x0546
		"11000100",	-- 0x0547
		"00010001",	-- 0x0548
		"01011110",	-- 0x0549
		"11111100",	-- 0x054A
		"00000001",	-- 0x054B
		"00001010",	-- 0x054C
		"00000000",	-- 0x054D
		"11101101",	-- 0x054E
		"10110000",	-- 0x054F
		"11001101",	-- 0x0550
		"01000001",	-- 0x0551
		"11000100",	-- 0x0552
		"00111010",	-- 0x0553
		"01101000",	-- 0x0554
		"11111100",	-- 0x0555
		"11111110",	-- 0x0556
		"00000111",	-- 0x0557
		"00100000",	-- 0x0558
		"01001010",	-- 0x0559
		"00111010",	-- 0x055A
		"01101001",	-- 0x055B
		"11111100",	-- 0x055C
		"11100110",	-- 0x055D
		"11000000",	-- 0x055E
		"00100000",	-- 0x055F
		"01000011",	-- 0x0560
		"00100001",	-- 0x0561
		"11101100",	-- 0x0562
		"11000100",	-- 0x0563
		"00010001",	-- 0x0564
		"01011110",	-- 0x0565
		"11111100",	-- 0x0566
		"00000001",	-- 0x0567
		"00000100",	-- 0x0568
		"00000000",	-- 0x0569
		"11101101",	-- 0x056A
		"10110000",	-- 0x056B
		"11001101",	-- 0x056C
		"00001010",	-- 0x056D
		"11000101",	-- 0x056E
		"00100001",	-- 0x056F
		"11110000",	-- 0x0570
		"11000100",	-- 0x0571
		"00001110",	-- 0x0572
		"11111111",	-- 0x0573
		"00000110",	-- 0x0574
		"00010000",	-- 0x0575
		"11101101",	-- 0x0576
		"10110011",	-- 0x0577
		"00100001",	-- 0x0578
		"00000000",	-- 0x0579
		"11000101",	-- 0x057A
		"00010001",	-- 0x057B
		"01011110",	-- 0x057C
		"11111100",	-- 0x057D
		"00000001",	-- 0x057E
		"00001010",	-- 0x057F
		"00000000",	-- 0x0580
		"11101101",	-- 0x0581
		"10110000",	-- 0x0582
		"11001101",	-- 0x0583
		"01000001",	-- 0x0584
		"11000100",	-- 0x0585
		"00111010",	-- 0x0586
		"01101000",	-- 0x0587
		"11111100",	-- 0x0588
		"11111110",	-- 0x0589
		"00000111",	-- 0x058A
		"00100000",	-- 0x058B
		"00010111",	-- 0x058C
		"00111010",	-- 0x058D
		"01101001",	-- 0x058E
		"11111100",	-- 0x058F
		"11100110",	-- 0x0590
		"11000000",	-- 0x0591
		"00100000",	-- 0x0592
		"00010000",	-- 0x0593
		"11001101",	-- 0x0594
		"01001000",	-- 0x0595
		"11000011",	-- 0x0596
		"00111010",	-- 0x0597
		"01011011",	-- 0x0598
		"11111100",	-- 0x0599
		"11001011",	-- 0x059A
		"10000111",	-- 0x059B
		"00110010",	-- 0x059C
		"01011011",	-- 0x059D
		"11111100",	-- 0x059E
		"11000001",	-- 0x059F
		"11000011",	-- 0x05A0
		"10000000",	-- 0x05A1
		"10011111",	-- 0x05A2
		"11100001",	-- 0x05A3
		"11000001",	-- 0x05A4
		"00010000",	-- 0x05A5
		"10010001",	-- 0x05A6
		"11011011",	-- 0x05A7
		"11101100",	-- 0x05A8
		"11101110",	-- 0x05A9
		"00000001",	-- 0x05AA
		"11010011",	-- 0x05AB
		"11101100",	-- 0x05AC
		"11000011",	-- 0x05AD
		"11111001",	-- 0x05AE
		"11000000",	-- 0x05AF
		"11110101",	-- 0x05B0
		"00111110",	-- 0x05B1
		"10100011",	-- 0x05B2
		"11010011",	-- 0x05B3
		"11111111",	-- 0x05B4
		"11110001",	-- 0x05B5
		"11111011",	-- 0x05B6
		"11101101",	-- 0x05B7
		"01001101",	-- 0x05B8
		"00111010",	-- 0x05B9
		"01011010",	-- 0x05BA
		"11111100",	-- 0x05BB
		"10110111",	-- 0x05BC
		"00101000",	-- 0x05BD
		"00000010",	-- 0x05BE
		"00111110",	-- 0x05BF
		"11111111",	-- 0x05C0
		"11111110",	-- 0x05C1
		"11111111",	-- 0x05C2
		"11001001",	-- 0x05C3
		"00000000",	-- 0x05C4
		"11110101",	-- 0x05C5
		"11000101",	-- 0x05C6
		"11010101",	-- 0x05C7
		"11100101",	-- 0x05C8
		"11001101",	-- 0x05C9
		"11000110",	-- 0x05CA
		"11000111",	-- 0x05CB
		"11100001",	-- 0x05CC
		"11010001",	-- 0x05CD
		"11000001",	-- 0x05CE
		"11110001",	-- 0x05CF
		"11001001",	-- 0x05D0
		"11110101",	-- 0x05D1
		"11000101",	-- 0x05D2
		"11010101",	-- 0x05D3
		"11100101",	-- 0x05D4
		"11001101",	-- 0x05D5
		"11111011",	-- 0x05D6
		"11000101",	-- 0x05D7
		"11001101",	-- 0x05D8
		"01010111",	-- 0x05D9
		"11001000",	-- 0x05DA
		"00111110",	-- 0x05DB
		"00011011",	-- 0x05DC
		"00110010",	-- 0x05DD
		"00100110",	-- 0x05DE
		"11111100",	-- 0x05DF
		"00011000",	-- 0x05E0
		"11101010",	-- 0x05E1
		"00001000",	-- 0x05E2
		"00010110",	-- 0x05E3
		"00101100",	-- 0x05E4
		"10000101",	-- 0x05E5
		"00010101",	-- 0x05E6
		"00000101",	-- 0x05E7
		"00000010",	-- 0x05E8
		"00001000",	-- 0x05E9
		"01111101",	-- 0x05EA
		"00001000",	-- 0x05EB
		"00010110",	-- 0x05EC
		"00101100",	-- 0x05ED
		"10000101",	-- 0x05EE
		"00000101",	-- 0x05EF
		"00000001",	-- 0x05F0
		"00101111",	-- 0x05F1
		"00001000",	-- 0x05F2
		"11000001",	-- 0x05F3
		"00000110",	-- 0x05F4
		"10000000",	-- 0x05F5
		"00010000",	-- 0x05F6
		"00000000",	-- 0x05F7
		"00000000",	-- 0x05F8
		"00000000",	-- 0x05F9
		"00000000",	-- 0x05FA
		"10101111",	-- 0x05FB
		"00110010",	-- 0x05FC
		"00001001",	-- 0x05FD
		"11111100",	-- 0x05FE
		"00110010",	-- 0x05FF
		"00001001",	-- 0x0600
		"11111100",	-- 0x0601
		"00110010",	-- 0x0602
		"00010101",	-- 0x0603
		"11111100",	-- 0x0604
		"00111100",	-- 0x0605
		"00110010",	-- 0x0606
		"00000000",	-- 0x0607
		"11111100",	-- 0x0608
		"00110010",	-- 0x0609
		"00010110",	-- 0x060A
		"11111100",	-- 0x060B
		"00110010",	-- 0x060C
		"00011100",	-- 0x060D
		"11111100",	-- 0x060E
		"00110010",	-- 0x060F
		"00000001",	-- 0x0610
		"11111100",	-- 0x0611
		"00111110",	-- 0x0612
		"00000000",	-- 0x0613
		"11010011",	-- 0x0614
		"01110001",	-- 0x0615
		"00001110",	-- 0x0616
		"01110000",	-- 0x0617
		"00100001",	-- 0x0618
		"11100010",	-- 0x0619
		"11000101",	-- 0x061A
		"11011011",	-- 0x061B
		"11100111",	-- 0x061C
		"11001011",	-- 0x061D
		"01101111",	-- 0x061E
		"00101000",	-- 0x061F
		"00000011",	-- 0x0620
		"00100001",	-- 0x0621
		"11101011",	-- 0x0622
		"11000101",	-- 0x0623
		"01000110",	-- 0x0624
		"00100011",	-- 0x0625
		"11101101",	-- 0x0626
		"10110011",	-- 0x0627
		"11001101",	-- 0x0628
		"11000100",	-- 0x0629
		"11000110",	-- 0x062A
		"00111110",	-- 0x062B
		"01101111",	-- 0x062C
		"11010011",	-- 0x062D
		"01110001",	-- 0x062E
		"00100001",	-- 0x062F
		"11110100",	-- 0x0630
		"11000101",	-- 0x0631
		"01000110",	-- 0x0632
		"00100011",	-- 0x0633
		"00111110",	-- 0x0634
		"01110010",	-- 0x0635
		"11010011",	-- 0x0636
		"01110001",	-- 0x0637
		"11101101",	-- 0x0638
		"10110011",	-- 0x0639
		"00111110",	-- 0x063A
		"01001010",	-- 0x063B
		"11010011",	-- 0x063C
		"01110001",	-- 0x063D
		"00111110",	-- 0x063E
		"11111111",	-- 0x063F
		"11101101",	-- 0x0640
		"01111001",	-- 0x0641
		"11101101",	-- 0x0642
		"01111001",	-- 0x0643
		"00111110",	-- 0x0644
		"01000111",	-- 0x0645
		"11010011",	-- 0x0646
		"01110001",	-- 0x0647
		"00111110",	-- 0x0648
		"00101110",	-- 0x0649
		"11101101",	-- 0x064A
		"01111001",	-- 0x064B
		"00100001",	-- 0x064C
		"00000000",	-- 0x064D
		"00000000",	-- 0x064E
		"00100010",	-- 0x064F
		"00000101",	-- 0x0650
		"11111100",	-- 0x0651
		"11001101",	-- 0x0652
		"10110100",	-- 0x0653
		"11000110",	-- 0x0654
		"00010001",	-- 0x0655
		"00000111",	-- 0x0656
		"00000001",	-- 0x0657
		"00100001",	-- 0x0658
		"01000010",	-- 0x0659
		"00101111",	-- 0x065A
		"11101101",	-- 0x065B
		"01001011",	-- 0x065C
		"00000101",	-- 0x065D
		"11111100",	-- 0x065E
		"00001001",	-- 0x065F
		"00100010",	-- 0x0660
		"00000010",	-- 0x0661
		"11111100",	-- 0x0662
		"10101111",	-- 0x0663
		"00110010",	-- 0x0664
		"00000100",	-- 0x0665
		"11111100",	-- 0x0666
		"11001101",	-- 0x0667
		"01111111",	-- 0x0668
		"11000111",	-- 0x0669
		"00111110",	-- 0x066A
		"00110000",	-- 0x066B
		"11010011",	-- 0x066C
		"01110001",	-- 0x066D
		"11001101",	-- 0x066E
		"11000100",	-- 0x066F
		"11000110",	-- 0x0670
		"00111110",	-- 0x0671
		"01001100",	-- 0x0672
		"11010011",	-- 0x0673
		"01110001",	-- 0x0674
		"00111110",	-- 0x0675
		"00010010",	-- 0x0676
		"11101101",	-- 0x0677
		"01111001",	-- 0x0678
		"11101101",	-- 0x0679
		"01011001",	-- 0x067A
		"11101101",	-- 0x067B
		"01010001",	-- 0x067C
		"00100001",	-- 0x067D
		"11100000",	-- 0x067E
		"00000010",	-- 0x067F
		"11101101",	-- 0x0680
		"01101001",	-- 0x0681
		"11101101",	-- 0x0682
		"01100001",	-- 0x0683
		"11101101",	-- 0x0684
		"01101001",	-- 0x0685
		"11101101",	-- 0x0686
		"01100001",	-- 0x0687
		"11001101",	-- 0x0688
		"11000100",	-- 0x0689
		"11000110",	-- 0x068A
		"00111110",	-- 0x068B
		"01000110",	-- 0x068C
		"11010011",	-- 0x068D
		"01110001",	-- 0x068E
		"10101111",	-- 0x068F
		"11101101",	-- 0x0690
		"01111001",	-- 0x0691
		"00111110",	-- 0x0692
		"01111000",	-- 0x0693
		"11010011",	-- 0x0694
		"01110001",	-- 0x0695
		"00000110",	-- 0x0696
		"00001000",	-- 0x0697
		"00111110",	-- 0x0698
		"00000000",	-- 0x0699
		"11101101",	-- 0x069A
		"01111001",	-- 0x069B
		"00010000",	-- 0x069C
		"11111100",	-- 0x069D
		"00100001",	-- 0x069E
		"01101000",	-- 0x069F
		"00001101",	-- 0x06A0
		"00001110",	-- 0x06A1
		"01110001",	-- 0x06A2
		"11101101",	-- 0x06A3
		"01101001",	-- 0x06A4
		"11101101",	-- 0x06A5
		"01100001",	-- 0x06A6
		"00111110",	-- 0x06A7
		"00000001",	-- 0x06A8
		"00110010",	-- 0x06A9
		"00000000",	-- 0x06AA
		"11111100",	-- 0x06AB
		"00111110",	-- 0x06AC
		"00000001",	-- 0x06AD
		"00110010",	-- 0x06AE
		"00000001",	-- 0x06AF
		"11111100",	-- 0x06B0
		"11000011",	-- 0x06B1
		"00101101",	-- 0x06B2
		"11000111",	-- 0x06B3
		"11001101",	-- 0x06B4
		"11000100",	-- 0x06B5
		"11000110",	-- 0x06B6
		"00111110",	-- 0x06B7
		"01110000",	-- 0x06B8
		"00100001",	-- 0x06B9
		"00000101",	-- 0x06BA
		"11111100",	-- 0x06BB
		"11010011",	-- 0x06BC
		"01110001",	-- 0x06BD
		"00000001",	-- 0x06BE
		"01110000",	-- 0x06BF
		"00000010",	-- 0x06C0
		"11101101",	-- 0x06C1
		"10110011",	-- 0x06C2
		"11001001",	-- 0x06C3
		"11011011",	-- 0x06C4
		"01110000",	-- 0x06C5
		"11001011",	-- 0x06C6
		"01010111",	-- 0x06C7
		"11000000",	-- 0x06C8
		"00011000",	-- 0x06C9
		"11111001",	-- 0x06CA
		"11011011",	-- 0x06CB
		"01110000",	-- 0x06CC
		"11001011",	-- 0x06CD
		"01001111",	-- 0x06CE
		"11001000",	-- 0x06CF
		"00011000",	-- 0x06D0
		"11111001",	-- 0x06D1
		"11011011",	-- 0x06D2
		"01110000",	-- 0x06D3
		"11001011",	-- 0x06D4
		"01000111",	-- 0x06D5
		"11001001",	-- 0x06D6
		"00010110",	-- 0x06D7
		"00000001",	-- 0x06D8
		"00011110",	-- 0x06D9
		"00001001",	-- 0x06DA
		"11001101",	-- 0x06DB
		"11000100",	-- 0x06DC
		"11000110",	-- 0x06DD
		"00111110",	-- 0x06DE
		"01000110",	-- 0x06DF
		"11010011",	-- 0x06E0
		"01110001",	-- 0x06E1
		"00111110",	-- 0x06E2
		"00000001",	-- 0x06E3
		"00111101",	-- 0x06E4
		"11010011",	-- 0x06E5
		"01110000",	-- 0x06E6
		"00111110",	-- 0x06E7
		"01001100",	-- 0x06E8
		"11010011",	-- 0x06E9
		"01110001",	-- 0x06EA
		"00001110",	-- 0x06EB
		"01110000",	-- 0x06EC
		"00111110",	-- 0x06ED
		"00010010",	-- 0x06EE
		"11101101",	-- 0x06EF
		"01111001",	-- 0x06F0
		"10101111",	-- 0x06F1
		"11101101",	-- 0x06F2
		"01010001",	-- 0x06F3
		"11101101",	-- 0x06F4
		"01111001",	-- 0x06F5
		"11101101",	-- 0x06F6
		"01011001",	-- 0x06F7
		"11101101",	-- 0x06F8
		"01111001",	-- 0x06F9
		"11101101",	-- 0x06FA
		"01011001",	-- 0x06FB
		"11101101",	-- 0x06FC
		"01111001",	-- 0x06FD
		"11001101",	-- 0x06FE
		"11000100",	-- 0x06FF
		"11000110",	-- 0x0700
		"00111110",	-- 0x0701
		"01111000",	-- 0x0702
		"11010011",	-- 0x0703
		"01110001",	-- 0x0704
		"00000110",	-- 0x0705
		"00001000",	-- 0x0706
		"00111110",	-- 0x0707
		"11111111",	-- 0x0708
		"11101101",	-- 0x0709
		"01111001",	-- 0x070A
		"00010000",	-- 0x070B
		"11111100",	-- 0x070C
		"11001101",	-- 0x070D
		"11001011",	-- 0x070E
		"11000110",	-- 0x070F
		"00111110",	-- 0x0710
		"00110001",	-- 0x0711
		"11010011",	-- 0x0712
		"01110001",	-- 0x0713
		"00111110",	-- 0x0714
		"01101000",	-- 0x0715
		"11010011",	-- 0x0716
		"01110001",	-- 0x0717
		"11001001",	-- 0x0718
		"00100001",	-- 0x0719
		"00000000",	-- 0x071A
		"00000000",	-- 0x071B
		"00111110",	-- 0x071C
		"00010001",	-- 0x071D
		"11001011",	-- 0x071E
		"00011000",	-- 0x071F
		"11001011",	-- 0x0720
		"00011001",	-- 0x0721
		"00111101",	-- 0x0722
		"11001000",	-- 0x0723
		"00110000",	-- 0x0724
		"00000001",	-- 0x0725
		"00011001",	-- 0x0726
		"11001011",	-- 0x0727
		"00011100",	-- 0x0728
		"11001011",	-- 0x0729
		"00011101",	-- 0x072A
		"00011000",	-- 0x072B
		"11110001",	-- 0x072C
		"00010001",	-- 0x072D
		"00001011",	-- 0x072E
		"00000000",	-- 0x072F
		"00000001",	-- 0x0730
		"00101110",	-- 0x0731
		"00000000",	-- 0x0732
		"11001101",	-- 0x0733
		"00011001",	-- 0x0734
		"11000111",	-- 0x0735
		"11101101",	-- 0x0736
		"01011011",	-- 0x0737
		"00000000",	-- 0x0738
		"11111100",	-- 0x0739
		"00010110",	-- 0x073A
		"00000000",	-- 0x073B
		"11001101",	-- 0x073C
		"00011001",	-- 0x073D
		"11000111",	-- 0x073E
		"01100000",	-- 0x073F
		"01101001",	-- 0x0740
		"00000001",	-- 0x0741
		"00101110",	-- 0x0742
		"00000000",	-- 0x0743
		"10100111",	-- 0x0744
		"11101101",	-- 0x0745
		"01000010",	-- 0x0746
		"11101101",	-- 0x0747
		"01001011",	-- 0x0748
		"00000101",	-- 0x0749
		"11111100",	-- 0x074A
		"00001001",	-- 0x074B
		"00100010",	-- 0x074C
		"00000111",	-- 0x074D
		"11111100",	-- 0x074E
		"10101111",	-- 0x074F
		"00011110",	-- 0x0750
		"00001001",	-- 0x0751
		"01010111",	-- 0x0752
		"11101101",	-- 0x0753
		"01001011",	-- 0x0754
		"00000001",	-- 0x0755
		"11111100",	-- 0x0756
		"01000111",	-- 0x0757
		"11001101",	-- 0x0758
		"00011001",	-- 0x0759
		"11000111",	-- 0x075A
		"01100000",	-- 0x075B
		"01101001",	-- 0x075C
		"10101111",	-- 0x075D
		"10101111",	-- 0x075E
		"11101101",	-- 0x075F
		"01010010",	-- 0x0760
		"00100010",	-- 0x0761
		"00011010",	-- 0x0762
		"11111100",	-- 0x0763
		"00000110",	-- 0x0764
		"00000100",	-- 0x0765
		"11001011",	-- 0x0766
		"00111100",	-- 0x0767
		"11001011",	-- 0x0768
		"00011101",	-- 0x0769
		"11001011",	-- 0x076A
		"00011111",	-- 0x076B
		"00010000",	-- 0x076C
		"11111000",	-- 0x076D
		"00110010",	-- 0x076E
		"00000100",	-- 0x076F
		"11111100",	-- 0x0770
		"00110010",	-- 0x0771
		"00011001",	-- 0x0772
		"11111100",	-- 0x0773
		"11101101",	-- 0x0774
		"01011011",	-- 0x0775
		"00000111",	-- 0x0776
		"11111100",	-- 0x0777
		"00011001",	-- 0x0778
		"00100010",	-- 0x0779
		"00000010",	-- 0x077A
		"11111100",	-- 0x077B
		"00100010",	-- 0x077C
		"00010111",	-- 0x077D
		"11111100",	-- 0x077E
		"11001101",	-- 0x077F
		"11000100",	-- 0x0780
		"11000110",	-- 0x0781
		"00111110",	-- 0x0782
		"01001001",	-- 0x0783
		"00100001",	-- 0x0784
		"00000010",	-- 0x0785
		"11111100",	-- 0x0786
		"11001101",	-- 0x0787
		"10111100",	-- 0x0788
		"11000110",	-- 0x0789
		"00111010",	-- 0x078A
		"00000100",	-- 0x078B
		"11111100",	-- 0x078C
		"11100110",	-- 0x078D
		"11110000",	-- 0x078E
		"11101101",	-- 0x078F
		"01111001",	-- 0x0790
		"11001001",	-- 0x0791
		"01111001",	-- 0x0792
		"00100001",	-- 0x0793
		"10111010",	-- 0x0794
		"11000111",	-- 0x0795
		"00000001",	-- 0x0796
		"00000100",	-- 0x0797
		"00000000",	-- 0x0798
		"11101101",	-- 0x0799
		"10110001",	-- 0x079A
		"11000000",	-- 0x079B
		"11000101",	-- 0x079C
		"11001101",	-- 0x079D
		"01101000",	-- 0x079E
		"11001000",	-- 0x079F
		"11001101",	-- 0x07A0
		"01111111",	-- 0x07A1
		"11000111",	-- 0x07A2
		"11000001",	-- 0x07A3
		"00100001",	-- 0x07A4
		"10111110",	-- 0x07A5
		"11000111",	-- 0x07A6
		"11001101",	-- 0x07A7
		"10110011",	-- 0x07A8
		"11000111",	-- 0x07A9
		"00101010",	-- 0x07AA
		"00011010",	-- 0x07AB
		"11111100",	-- 0x07AC
		"11001101",	-- 0x07AD
		"01100001",	-- 0x07AE
		"11000111",	-- 0x07AF
		"11000011",	-- 0x07B0
		"01010111",	-- 0x07B1
		"11001000",	-- 0x07B2
		"00001001",	-- 0x07B3
		"00001001",	-- 0x07B4
		"01001110",	-- 0x07B5
		"00100011",	-- 0x07B6
		"01100110",	-- 0x07B7
		"01101001",	-- 0x07B8
		"11101001",	-- 0x07B9
		"00001010",	-- 0x07BA
		"00001101",	-- 0x07BB
		"00001100",	-- 0x07BC
		"00000111",	-- 0x07BD
		"00010111",	-- 0x07BE
		"11001001",	-- 0x07BF
		"01010101",	-- 0x07C0
		"11000110",	-- 0x07C1
		"11111110",	-- 0x07C2
		"11001000",	-- 0x07C3
		"00000101",	-- 0x07C4
		"11001001",	-- 0x07C5
		"01111001",	-- 0x07C6
		"11111110",	-- 0x07C7
		"00100000",	-- 0x07C8
		"11011010",	-- 0x07C9
		"10010010",	-- 0x07CA
		"11000111",	-- 0x07CB
		"11001011",	-- 0x07CC
		"10111001",	-- 0x07CD
		"11001101",	-- 0x07CE
		"11010100",	-- 0x07CF
		"11000111",	-- 0x07D0
		"11000011",	-- 0x07D1
		"01000010",	-- 0x07D2
		"11001000",	-- 0x07D3
		"00101010",	-- 0x07D4
		"00110110",	-- 0x07D5
		"11001001",	-- 0x07D6
		"00000110",	-- 0x07D7
		"00000000",	-- 0x07D8
		"00001001",	-- 0x07D9
		"00001001",	-- 0x07DA
		"01011110",	-- 0x07DB
		"00100011",	-- 0x07DC
		"01100110",	-- 0x07DD
		"01101011",	-- 0x07DE
		"00000001",	-- 0x07DF
		"00001011",	-- 0x07E0
		"00000000",	-- 0x07E1
		"00010001",	-- 0x07E2
		"00001010",	-- 0x07E3
		"11111100",	-- 0x07E4
		"11101101",	-- 0x07E5
		"10110000",	-- 0x07E6
		"11001101",	-- 0x07E7
		"11000100",	-- 0x07E8
		"11000110",	-- 0x07E9
		"00111110",	-- 0x07EA
		"01000110",	-- 0x07EB
		"11010011",	-- 0x07EC
		"01110001",	-- 0x07ED
		"00111110",	-- 0x07EE
		"00000001",	-- 0x07EF
		"00111101",	-- 0x07F0
		"11010011",	-- 0x07F1
		"01110000",	-- 0x07F2
		"00111110",	-- 0x07F3
		"00110000",	-- 0x07F4
		"11010011",	-- 0x07F5
		"01110001",	-- 0x07F6
		"00011110",	-- 0x07F7
		"00001001",	-- 0x07F8
		"00111110",	-- 0x07F9
		"00010010",	-- 0x07FA
		"01010111",	-- 0x07FB
		"11001101",	-- 0x07FC
		"01111111",	-- 0x07FD
		"11000111",	-- 0x07FE
		"00000001",	-- 0x07FF
		"11110011",	-- 0x0800
		"11000011",	-- 0x0801
		"00010011",	-- 0x0802
		"11000000",	-- 0x0803
		"11000011",	-- 0x0804
		"00011010",	-- 0x0805
		"11000100",	-- 0x0806
		"11000011",	-- 0x0807
		"11100110",	-- 0x0808
		"11111100",	-- 0x0809
		"11000011",	-- 0x080A
		"00110100",	-- 0x080B
		"11000100",	-- 0x080C
		"11000011",	-- 0x080D
		"00111110",	-- 0x080E
		"11000100",	-- 0x080F
		"11000011",	-- 0x0810
		"10010101",	-- 0x0811
		"11000000",	-- 0x0812
		"00111110",	-- 0x0813
		"11001111",	-- 0x0814
		"11010011",	-- 0x0815
		"11101110",	-- 0x0816
		"00111110",	-- 0x0817
		"10000000",	-- 0x0818
		"11010011",	-- 0x0819
		"11101110",	-- 0x081A
		"00111110",	-- 0x081B
		"01000000",	-- 0x081C
		"11010011",	-- 0x081D
		"11101100",	-- 0x081E
		"11000011",	-- 0x081F
		"01001111",	-- 0x0820
		"11000000",	-- 0x0821
		"11000011",	-- 0x0822
		"10111001",	-- 0x0823
		"11000101",	-- 0x0824
		"11011011",	-- 0x0825
		"11111110",	-- 0x0826
		"01111110",	-- 0x0827
		"11010011",	-- 0x0828
		"11111110",	-- 0x0829
		"11001001",	-- 0x082A
		"11011011",	-- 0x082B
		"11111110",	-- 0x082C
		"01110001",	-- 0x082D
		"11010011",	-- 0x082E
		"11111110",	-- 0x082F
		"11001001",	-- 0x0830
		"11000011",	-- 0x0831
		"10111110",	-- 0x0832
		"11000011",	-- 0x0833
		"01001111",	-- 0x0834
		"11000011",	-- 0x0835
		"11000101",	-- 0x0836
		"11000101",	-- 0x0837
		"11000011",	-- 0x0838
		"00011101",	-- 0x0839
		"11000100",	-- 0x083A
		"00001101",	-- 0x083B
		"01001101",	-- 0x083C
		"01001111",	-- 0x083D
		"01001110",	-- 0x083E
		"01001001",	-- 0x083F
		"00100000",	-- 0x0840
		"01001101",	-- 0x0841
		"01010000",	-- 0x0842
		"01000011",	-- 0x0843
		"00100000",	-- 0x0844
		"01010110",	-- 0x0845
		"00101110",	-- 0x0846
		"00110000",	-- 0x0847
		"00110001",	-- 0x0848
		"00001101",	-- 0x0849
		"00001101",	-- 0x084A
		"01001001",	-- 0x084B
		"01001110",	-- 0x084C
		"01001001",	-- 0x084D
		"01010100",	-- 0x084E
		"00100001",	-- 0x084F
		"01011010",	-- 0x0850
		"11111100",	-- 0x0851
		"00000110",	-- 0x0852
		"10000010",	-- 0x0853
		"10101111",	-- 0x0854
		"01110111",	-- 0x0855
		"00100011",	-- 0x0856
		"00010000",	-- 0x0857
		"11111011",	-- 0x0858
		"00110001",	-- 0x0859
		"11011100",	-- 0x085A
		"11111100",	-- 0x085B
		"11001101",	-- 0x085C
		"11101111",	-- 0x085D
		"11000011",	-- 0x085E
		"00100001",	-- 0x085F
		"00100010",	-- 0x0860
		"11000000",	-- 0x0861
		"00010001",	-- 0x0862
		"11100110",	-- 0x0863
		"11111100",	-- 0x0864
		"00000001",	-- 0x0865
		"00011001",	-- 0x0866
		"00000000",	-- 0x0867
		"11101101",	-- 0x0868
		"10110000",	-- 0x0869
		"00100001",	-- 0x086A
		"10110000",	-- 0x086B
		"11000101",	-- 0x086C
		"00010001",	-- 0x086D
		"11011100",	-- 0x086E
		"11111100",	-- 0x086F
		"00000001",	-- 0x0870
		"00001001",	-- 0x0871
		"00000000",	-- 0x0872
		"11101101",	-- 0x0873
		"10110000",	-- 0x0874
		"00100001",	-- 0x0875
		"01001010",	-- 0x0876
		"11000000",	-- 0x0877
		"00000110",	-- 0x0878
		"00000101",	-- 0x0879
		"11001101",	-- 0x087A
		"00111100",	-- 0x087B
		"11000011",	-- 0x087C
		"00111110",	-- 0x087D
		"11000011",	-- 0x087E
		"00100001",	-- 0x087F
		"10010101",	-- 0x0880
		"11000000",	-- 0x0881
		"00110010",	-- 0x0882
		"00111000",	-- 0x0883
		"00000000",	-- 0x0884
		"00100010",	-- 0x0885
		"00111001",	-- 0x0886
		"00000000",	-- 0x0887
		"00111110",	-- 0x0888
		"10000001",	-- 0x0889
		"00110010",	-- 0x088A
		"01011011",	-- 0x088B
		"11111100",	-- 0x088C
		"00100001",	-- 0x088D
		"00000000",	-- 0x088E
		"00000000",	-- 0x088F
		"00111110",	-- 0x0890
		"11111101",	-- 0x0891
		"11101101",	-- 0x0892
		"01000111",	-- 0x0893
		"11100101",	-- 0x0894
		"11110011",	-- 0x0895
		"11101101",	-- 0x0896
		"01011110",	-- 0x0897
		"00100010",	-- 0x0898
		"01001110",	-- 0x0899
		"11111100",	-- 0x089A
		"11100001",	-- 0x089B
		"00100010",	-- 0x089C
		"01010110",	-- 0x089D
		"11111100",	-- 0x089E
		"11101101",	-- 0x089F
		"01110011",	-- 0x08A0
		"01011000",	-- 0x08A1
		"11111100",	-- 0x08A2
		"00110001",	-- 0x08A3
		"01010110",	-- 0x08A4
		"11111100",	-- 0x08A5
		"11110101",	-- 0x08A6
		"11000101",	-- 0x08A7
		"11010101",	-- 0x08A8
		"00001000",	-- 0x08A9
		"11011001",	-- 0x08AA
		"00111011",	-- 0x08AB
		"00111011",	-- 0x08AC
		"11110101",	-- 0x08AD
		"11000101",	-- 0x08AE
		"11010101",	-- 0x08AF
		"11100101",	-- 0x08B0
		"11011101",	-- 0x08B1
		"11100101",	-- 0x08B2
		"11111101",	-- 0x08B3
		"11100101",	-- 0x08B4
		"11101101",	-- 0x08B5
		"01010111",	-- 0x08B6
		"11110101",	-- 0x08B7
		"00111110",	-- 0x08B8
		"11111101",	-- 0x08B9
		"11101101",	-- 0x08BA
		"01000111",	-- 0x08BB
		"00111010",	-- 0x08BC
		"01011011",	-- 0x08BD
		"11111100",	-- 0x08BE
		"11001011",	-- 0x08BF
		"11000111",	-- 0x08C0
		"00110010",	-- 0x08C1
		"01011011",	-- 0x08C2
		"11111100",	-- 0x08C3
		"00110001",	-- 0x08C4
		"10011110",	-- 0x08C5
		"11111100",	-- 0x08C6
		"11111011",	-- 0x08C7
		"00100001",	-- 0x08C8
		"00111011",	-- 0x08C9
		"11000000",	-- 0x08CA
		"00000110",	-- 0x08CB
		"00001111",	-- 0x08CC
		"11001101",	-- 0x08CD
		"00111100",	-- 0x08CE
		"11000011",	-- 0x08CF
		"00100001",	-- 0x08D0
		"01011011",	-- 0x08D1
		"11111100",	-- 0x08D2
		"11001011",	-- 0x08D3
		"01111110",	-- 0x08D4
		"11001011",	-- 0x08D5
		"10111110",	-- 0x08D6
		"11000010",	-- 0x08D7
		"00110110",	-- 0x08D8
		"11000101",	-- 0x08D9
		"00111110",	-- 0x08DA
		"00111010",	-- 0x08DB
		"11001101",	-- 0x08DC
		"00110111",	-- 0x08DD
		"11000001",	-- 0x08DE
		"11001101",	-- 0x08DF
		"00011111",	-- 0x08E0
		"11000001",	-- 0x08E1
		"11001101",	-- 0x08E2
		"11100000",	-- 0x08E3
		"11000011",	-- 0x08E4
		"00100001",	-- 0x08E5
		"00000100",	-- 0x08E6
		"11000001",	-- 0x08E7
		"00000001",	-- 0x08E8
		"00001001",	-- 0x08E9
		"00000000",	-- 0x08EA
		"11101101",	-- 0x08EB
		"10110001",	-- 0x08EC
		"00100000",	-- 0x08ED
		"00001010",	-- 0x08EE
		"00100001",	-- 0x08EF
		"00001101",	-- 0x08F0
		"11000001",	-- 0x08F1
		"00001001",	-- 0x08F2
		"00001001",	-- 0x08F3
		"01111110",	-- 0x08F4
		"00100011",	-- 0x08F5
		"01100110",	-- 0x08F6
		"01101111",	-- 0x08F7
		"11101001",	-- 0x08F8
		"00110001",	-- 0x08F9
		"10011110",	-- 0x08FA
		"11111100",	-- 0x08FB
		"00111110",	-- 0x08FC
		"00111111",	-- 0x08FD
		"11001101",	-- 0x08FE
		"00110111",	-- 0x08FF
		"11000001",	-- 0x0900
		"11000011",	-- 0x0901
		"01100001",	-- 0x0902
		"11000010",	-- 0x0903
		"01001100",	-- 0x0904
		"01001001",	-- 0x0905
		"01001111",	-- 0x0906
		"01000111",	-- 0x0907
		"01000100",	-- 0x0908
		"01000110",	-- 0x0909
		"01001101",	-- 0x090A
		"01010011",	-- 0x090B
		"01011000",	-- 0x090C
		"11001110",	-- 0x090D
		"11000010",	-- 0x090E
		"10100000",	-- 0x090F
		"11000010",	-- 0x0910
		"10000110",	-- 0x0911
		"11000010",	-- 0x0912
		"01110111",	-- 0x0913
		"11000010",	-- 0x0914
		"00001011",	-- 0x0915
		"11000010",	-- 0x0916
		"10001101",	-- 0x0917
		"11000011",	-- 0x0918
		"11010111",	-- 0x0919
		"11000011",	-- 0x091A
		"11001100",	-- 0x091B
		"11000011",	-- 0x091C
		"00110110",	-- 0x091D
		"11000101",	-- 0x091E
		"11000101",	-- 0x091F
		"11010101",	-- 0x0920
		"11001101",	-- 0x0921
		"01001110",	-- 0x0922
		"11000001",	-- 0x0923
		"11001101",	-- 0x0924
		"01000001",	-- 0x0925
		"11000001",	-- 0x0926
		"11010001",	-- 0x0927
		"11000001",	-- 0x0928
		"11001001",	-- 0x0929
		"00011010",	-- 0x092A
		"11110101",	-- 0x092B
		"00001111",	-- 0x092C
		"00001111",	-- 0x092D
		"00001111",	-- 0x092E
		"00001111",	-- 0x092F
		"11001101",	-- 0x0930
		"00110100",	-- 0x0931
		"11000001",	-- 0x0932
		"11110001",	-- 0x0933
		"11001101",	-- 0x0934
		"01010111",	-- 0x0935
		"11000001",	-- 0x0936
		"11110101",	-- 0x0937
		"11000101",	-- 0x0938
		"11010101",	-- 0x0939
		"11001101",	-- 0x093A
		"01000001",	-- 0x093B
		"11000001",	-- 0x093C
		"11010001",	-- 0x093D
		"11000001",	-- 0x093E
		"11110001",	-- 0x093F
		"11001001",	-- 0x0940
		"11001101",	-- 0x0941
		"00110100",	-- 0x0942
		"11000100",	-- 0x0943
		"11111110",	-- 0x0944
		"00001101",	-- 0x0945
		"11110101",	-- 0x0946
		"00111110",	-- 0x0947
		"00001010",	-- 0x0948
		"11001100",	-- 0x0949
		"00110100",	-- 0x094A
		"11000100",	-- 0x094B
		"11110001",	-- 0x094C
		"11001001",	-- 0x094D
		"11001101",	-- 0x094E
		"00011010",	-- 0x094F
		"11000100",	-- 0x0950
		"11111110",	-- 0x0951
		"00001101",	-- 0x0952
		"11000000",	-- 0x0953
		"11110101",	-- 0x0954
		"00011000",	-- 0x0955
		"11110010",	-- 0x0956
		"11100110",	-- 0x0957
		"00001111",	-- 0x0958
		"11000110",	-- 0x0959
		"00110000",	-- 0x095A
		"11111110",	-- 0x095B
		"00111010",	-- 0x095C
		"11111000",	-- 0x095D
		"11000110",	-- 0x095E
		"00000111",	-- 0x095F
		"11001001",	-- 0x0960
		"11010110",	-- 0x0961
		"00110000",	-- 0x0962
		"11111110",	-- 0x0963
		"00001010",	-- 0x0964
		"11111000",	-- 0x0965
		"11010110",	-- 0x0966
		"00000111",	-- 0x0967
		"11001001",	-- 0x0968
		"01111001",	-- 0x0969
		"11111110",	-- 0x096A
		"00110000",	-- 0x096B
		"00111111",	-- 0x096C
		"11010000",	-- 0x096D
		"11111110",	-- 0x096E
		"00111010",	-- 0x096F
		"11011000",	-- 0x0970
		"11111110",	-- 0x0971
		"01000001",	-- 0x0972
		"00111111",	-- 0x0973
		"11010000",	-- 0x0974
		"11111110",	-- 0x0975
		"01000111",	-- 0x0976
		"11001001",	-- 0x0977
		"11111110",	-- 0x0978
		"00110000",	-- 0x0979
		"00111111",	-- 0x097A
		"11010000",	-- 0x097B
		"11111110",	-- 0x097C
		"00111010",	-- 0x097D
		"11001001",	-- 0x097E
		"01111001",	-- 0x097F
		"11111110",	-- 0x0980
		"00101100",	-- 0x0981
		"00110111",	-- 0x0982
		"11001000",	-- 0x0983
		"11111110",	-- 0x0984
		"00100000",	-- 0x0985
		"00110111",	-- 0x0986
		"11001000",	-- 0x0987
		"11111110",	-- 0x0988
		"00001101",	-- 0x0989
		"00110111",	-- 0x098A
		"11001000",	-- 0x098B
		"00111111",	-- 0x098C
		"11001001",	-- 0x098D
		"11100101",	-- 0x098E
		"10110111",	-- 0x098F
		"11101101",	-- 0x0990
		"01010010",	-- 0x0991
		"00111111",	-- 0x0992
		"11100001",	-- 0x0993
		"11001001",	-- 0x0994
		"11100101",	-- 0x0995
		"00100001",	-- 0x0996
		"00000000",	-- 0x0997
		"00000000",	-- 0x0998
		"01011100",	-- 0x0999
		"11001101",	-- 0x099A
		"00011111",	-- 0x099B
		"11000001",	-- 0x099C
		"11001101",	-- 0x099D
		"11100000",	-- 0x099E
		"11000011",	-- 0x099F
		"01001111",	-- 0x09A0
		"11001101",	-- 0x09A1
		"01111111",	-- 0x09A2
		"11000001",	-- 0x09A3
		"00110000",	-- 0x09A4
		"00001001",	-- 0x09A5
		"01010001",	-- 0x09A6
		"11100101",	-- 0x09A7
		"11000001",	-- 0x09A8
		"11100001",	-- 0x09A9
		"01111011",	-- 0x09AA
		"10110111",	-- 0x09AB
		"11001000",	-- 0x09AC
		"00110111",	-- 0x09AD
		"11001001",	-- 0x09AE
		"11001101",	-- 0x09AF
		"01101001",	-- 0x09B0
		"11000001",	-- 0x09B1
		"11010010",	-- 0x09B2
		"11111001",	-- 0x09B3
		"11000000",	-- 0x09B4
		"01111001",	-- 0x09B5
		"11001101",	-- 0x09B6
		"01100001",	-- 0x09B7
		"11000001",	-- 0x09B8
		"00011110",	-- 0x09B9
		"11111111",	-- 0x09BA
		"00101001",	-- 0x09BB
		"00101001",	-- 0x09BC
		"00101001",	-- 0x09BD
		"00101001",	-- 0x09BE
		"00000110",	-- 0x09BF
		"00000000",	-- 0x09C0
		"01001111",	-- 0x09C1
		"00001001",	-- 0x09C2
		"00011000",	-- 0x09C3
		"11010101",	-- 0x09C4
		"01111100",	-- 0x09C5
		"11001101",	-- 0x09C6
		"00101011",	-- 0x09C7
		"11000001",	-- 0x09C8
		"01111101",	-- 0x09C9
		"11000011",	-- 0x09CA
		"00101011",	-- 0x09CB
		"11000001",	-- 0x09CC
		"00101110",	-- 0x09CD
		"00000011",	-- 0x09CE
		"01111001",	-- 0x09CF
		"11100110",	-- 0x09D0
		"00000011",	-- 0x09D1
		"01100111",	-- 0x09D2
		"11001101",	-- 0x09D3
		"10010101",	-- 0x09D4
		"11000001",	-- 0x09D5
		"11010010",	-- 0x09D6
		"11111001",	-- 0x09D7
		"11000000",	-- 0x09D8
		"11000101",	-- 0x09D9
		"00101101",	-- 0x09DA
		"00100101",	-- 0x09DB
		"01111010",	-- 0x09DC
		"00101000",	-- 0x09DD
		"00001010",	-- 0x09DE
		"11111110",	-- 0x09DF
		"00001101",	-- 0x09E0
		"11001010",	-- 0x09E1
		"11111001",	-- 0x09E2
		"11000000",	-- 0x09E3
		"00110010",	-- 0x09E4
		"01011100",	-- 0x09E5
		"11111100",	-- 0x09E6
		"00011000",	-- 0x09E7
		"11101010",	-- 0x09E8
		"11111110",	-- 0x09E9
		"00001101",	-- 0x09EA
		"11000010",	-- 0x09EB
		"11111001",	-- 0x09EC
		"11000000",	-- 0x09ED
		"00000001",	-- 0x09EE
		"11111111",	-- 0x09EF
		"11111111",	-- 0x09F0
		"01111101",	-- 0x09F1
		"10110111",	-- 0x09F2
		"00101000",	-- 0x09F3
		"00000100",	-- 0x09F4
		"11000101",	-- 0x09F5
		"00101101",	-- 0x09F6
		"00100000",	-- 0x09F7
		"11111100",	-- 0x09F8
		"11000001",	-- 0x09F9
		"11010001",	-- 0x09FA
		"11100001",	-- 0x09FB
		"11001101",	-- 0x09FC
		"10001110",	-- 0x09FD
		"11000001",	-- 0x09FE
		"00110000",	-- 0x09FF
		"00000000",	-- 0x0A00
		"11100011",	-- 0x0A01
		"11010101",	-- 0x0A02
		"11000101",	-- 0x0A03
		"11100101",	-- 0x0A04
		"00111101",	-- 0x0A05
		"11111000",	-- 0x0A06
		"11100001",	-- 0x0A07
		"11100011",	-- 0x0A08
		"00011000",	-- 0x0A09
		"11111010",	-- 0x0A0A
		"11001101",	-- 0x0A0B
		"01100111",	-- 0x0A0C
		"11000010",	-- 0x0A0D
		"11000101",	-- 0x0A0E
		"11000001",	-- 0x0A0F
		"00000110",	-- 0x0A10
		"00000000",	-- 0x0A11
		"11100101",	-- 0x0A12
		"11001101",	-- 0x0A13
		"11000101",	-- 0x0A14
		"11000001",	-- 0x0A15
		"10101111",	-- 0x0A16
		"10110000",	-- 0x0A17
		"11000100",	-- 0x0A18
		"01000100",	-- 0x0A19
		"11000011",	-- 0x0A1A
		"11001101",	-- 0x0A1B
		"01000100",	-- 0x0A1C
		"11000011",	-- 0x0A1D
		"11001101",	-- 0x0A1E
		"11101001",	-- 0x0A1F
		"11111100",	-- 0x0A20
		"00100000",	-- 0x0A21
		"00100000",	-- 0x0A22
		"11001101",	-- 0x0A23
		"00101011",	-- 0x0A24
		"11000001",	-- 0x0A25
		"11001101",	-- 0x0A26
		"10001110",	-- 0x0A27
		"11000001",	-- 0x0A28
		"00111000",	-- 0x0A29
		"00101010",	-- 0x0A2A
		"00100011",	-- 0x0A2B
		"01111101",	-- 0x0A2C
		"11100110",	-- 0x0A2D
		"00001111",	-- 0x0A2E
		"00100000",	-- 0x0A2F
		"11100101",	-- 0x0A30
		"11001101",	-- 0x0A31
		"01001000",	-- 0x0A32
		"11000011",	-- 0x0A33
		"00111010",	-- 0x0A34
		"01011100",	-- 0x0A35
		"11111100",	-- 0x0A36
		"11111110",	-- 0x0A37
		"00101100",	-- 0x0A38
		"00100000",	-- 0x0A39
		"11011000",	-- 0x0A3A
		"10101111",	-- 0x0A3B
		"10110000",	-- 0x0A3C
		"00100000",	-- 0x0A3D
		"11010000",	-- 0x0A3E
		"00000100",	-- 0x0A3F
		"11100001",	-- 0x0A40
		"00011000",	-- 0x0A41
		"11001111",	-- 0x0A42
		"11111110",	-- 0x0A43
		"00100000",	-- 0x0A44
		"00111000",	-- 0x0A45
		"00001001",	-- 0x0A46
		"11111110",	-- 0x0A47
		"01111111",	-- 0x0A48
		"00110000",	-- 0x0A49
		"00000101",	-- 0x0A4A
		"11001101",	-- 0x0A4B
		"00110111",	-- 0x0A4C
		"11000001",	-- 0x0A4D
		"00011000",	-- 0x0A4E
		"11010110",	-- 0x0A4F
		"11001101",	-- 0x0A50
		"01000100",	-- 0x0A51
		"11000011",	-- 0x0A52
		"00011000",	-- 0x0A53
		"11010001",	-- 0x0A54
		"00111010",	-- 0x0A55
		"01011100",	-- 0x0A56
		"11111100",	-- 0x0A57
		"11111110",	-- 0x0A58
		"00101100",	-- 0x0A59
		"00100000",	-- 0x0A5A
		"00000100",	-- 0x0A5B
		"10101111",	-- 0x0A5C
		"10110000",	-- 0x0A5D
		"00101000",	-- 0x0A5E
		"11010001",	-- 0x0A5F
		"11100001",	-- 0x0A60
		"11001101",	-- 0x0A61
		"01001000",	-- 0x0A62
		"11000011",	-- 0x0A63
		"11000011",	-- 0x0A64
		"11011010",	-- 0x0A65
		"11000000",	-- 0x0A66
		"00001110",	-- 0x0A67
		"00000010",	-- 0x0A68
		"11001101",	-- 0x0A69
		"11001101",	-- 0x0A6A
		"11000001",	-- 0x0A6B
		"11010001",	-- 0x0A6C
		"11100001",	-- 0x0A6D
		"11001001",	-- 0x0A6E
		"00001110",	-- 0x0A6F
		"00000011",	-- 0x0A70
		"11001101",	-- 0x0A71
		"11001101",	-- 0x0A72
		"11000001",	-- 0x0A73
		"11000001",	-- 0x0A74
		"00011000",	-- 0x0A75
		"11110101",	-- 0x0A76
		"11001101",	-- 0x0A77
		"01101111",	-- 0x0A78
		"11000010",	-- 0x0A79
		"11001101",	-- 0x0A7A
		"11101111",	-- 0x0A7B
		"11111100",	-- 0x0A7C
		"11001101",	-- 0x0A7D
		"10001110",	-- 0x0A7E
		"11000001",	-- 0x0A7F
		"11011010",	-- 0x0A80
		"11011010",	-- 0x0A81
		"11000000",	-- 0x0A82
		"00100011",	-- 0x0A83
		"00011000",	-- 0x0A84
		"11110100",	-- 0x0A85
		"11001101",	-- 0x0A86
		"01101111",	-- 0x0A87
		"11000010",	-- 0x0A88
		"11001101",	-- 0x0A89
		"11101001",	-- 0x0A8A
		"11111100",	-- 0x0A8B
		"11100101",	-- 0x0A8C
		"11000101",	-- 0x0A8D
		"01100000",	-- 0x0A8E
		"01101001",	-- 0x0A8F
		"01001111",	-- 0x0A90
		"11001101",	-- 0x0A91
		"11101111",	-- 0x0A92
		"11111100",	-- 0x0A93
		"11000001",	-- 0x0A94
		"11100001",	-- 0x0A95
		"00000011",	-- 0x0A96
		"11001101",	-- 0x0A97
		"10001110",	-- 0x0A98
		"11000001",	-- 0x0A99
		"00100011",	-- 0x0A9A
		"00100000",	-- 0x0A9B
		"11101100",	-- 0x0A9C
		"11000011",	-- 0x0A9D
		"11011010",	-- 0x0A9E
		"11000000",	-- 0x0A9F
		"11001101",	-- 0x0AA0
		"10010101",	-- 0x0AA1
		"11000001",	-- 0x0AA2
		"11000101",	-- 0x0AA3
		"11100001",	-- 0x0AA4
		"01111010",	-- 0x0AA5
		"11111110",	-- 0x0AA6
		"00001101",	-- 0x0AA7
		"11001010",	-- 0x0AA8
		"11011010",	-- 0x0AA9
		"11000000",	-- 0x0AAA
		"11001101",	-- 0x0AAB
		"11101001",	-- 0x0AAC
		"11111100",	-- 0x0AAD
		"11001101",	-- 0x0AAE
		"00101011",	-- 0x0AAF
		"11000001",	-- 0x0AB0
		"11001101",	-- 0x0AB1
		"10111100",	-- 0x0AB2
		"11000010",	-- 0x0AB3
		"00110000",	-- 0x0AB4
		"00000011",	-- 0x0AB5
		"11001101",	-- 0x0AB6
		"11101111",	-- 0x0AB7
		"11111100",	-- 0x0AB8
		"00100011",	-- 0x0AB9
		"00011000",	-- 0x0ABA
		"11101001",	-- 0x0ABB
		"00111110",	-- 0x0ABC
		"00101101",	-- 0x0ABD
		"11001101",	-- 0x0ABE
		"00110111",	-- 0x0ABF
		"11000001",	-- 0x0AC0
		"11000011",	-- 0x0AC1
		"10010101",	-- 0x0AC2
		"11000001",	-- 0x0AC3
		"00000110",	-- 0x0AC4
		"00000010",	-- 0x0AC5
		"11001101",	-- 0x0AC6
		"00111100",	-- 0x0AC7
		"11000011",	-- 0x0AC8
		"00111110",	-- 0x0AC9
		"00111101",	-- 0x0ACA
		"11000011",	-- 0x0ACB
		"00110111",	-- 0x0ACC
		"11000001",	-- 0x0ACD
		"11001101",	-- 0x0ACE
		"00011111",	-- 0x0ACF
		"11000001",	-- 0x0AD0
		"11001101",	-- 0x0AD1
		"11100000",	-- 0x0AD2
		"11000011",	-- 0x0AD3
		"11111110",	-- 0x0AD4
		"00001101",	-- 0x0AD5
		"00100001",	-- 0x0AD6
		"01001101",	-- 0x0AD7
		"11000011",	-- 0x0AD8
		"00010001",	-- 0x0AD9
		"01011001",	-- 0x0ADA
		"11111100",	-- 0x0ADB
		"00100000",	-- 0x0ADC
		"00000110",	-- 0x0ADD
		"11001101",	-- 0x0ADE
		"00011101",	-- 0x0ADF
		"11000011",	-- 0x0AE0
		"11000011",	-- 0x0AE1
		"11011010",	-- 0x0AE2
		"11000000",	-- 0x0AE3
		"11111110",	-- 0x0AE4
		"00100000",	-- 0x0AE5
		"00101000",	-- 0x0AE6
		"00000011",	-- 0x0AE7
		"11000011",	-- 0x0AE8
		"11111001",	-- 0x0AE9
		"11000000",	-- 0x0AEA
		"11001101",	-- 0x0AEB
		"11000100",	-- 0x0AEC
		"11000010",	-- 0x0AED
		"11001101",	-- 0x0AEE
		"00101010",	-- 0x0AEF
		"11000001",	-- 0x0AF0
		"11001011",	-- 0x0AF1
		"01000110",	-- 0x0AF2
		"00101000",	-- 0x0AF3
		"00000100",	-- 0x0AF4
		"00011011",	-- 0x0AF5
		"11001101",	-- 0x0AF6
		"00101010",	-- 0x0AF7
		"11000001",	-- 0x0AF8
		"11010101",	-- 0x0AF9
		"11001101",	-- 0x0AFA
		"10111100",	-- 0x0AFB
		"11000010",	-- 0x0AFC
		"01111010",	-- 0x0AFD
		"00110000",	-- 0x0AFE
		"00001111",	-- 0x0AFF
		"11010001",	-- 0x0B00
		"11110101",	-- 0x0B01
		"01111110",	-- 0x0B02
		"11101011",	-- 0x0B03
		"01110001",	-- 0x0B04
		"11001011",	-- 0x0B05
		"01000111",	-- 0x0B06
		"00101000",	-- 0x0B07
		"00000011",	-- 0x0B08
		"00100011",	-- 0x0B09
		"01110000",	-- 0x0B0A
		"00101011",	-- 0x0B0B
		"11110001",	-- 0x0B0C
		"11101011",	-- 0x0B0D
		"11010101",	-- 0x0B0E
		"11010001",	-- 0x0B0F
		"00011011",	-- 0x0B10
		"00100011",	-- 0x0B11
		"11111110",	-- 0x0B12
		"00001101",	-- 0x0B13
		"00101000",	-- 0x0B14
		"11001011",	-- 0x0B15
		"10101111",	-- 0x0B16
		"10110110",	-- 0x0B17
		"11001010",	-- 0x0B18
		"01100001",	-- 0x0B19
		"11000010",	-- 0x0B1A
		"00011000",	-- 0x0B1B
		"11001110",	-- 0x0B1C
		"01111110",	-- 0x0B1D
		"10110111",	-- 0x0B1E
		"11001010",	-- 0x0B1F
		"01001000",	-- 0x0B20
		"11000011",	-- 0x0B21
		"11001101",	-- 0x0B22
		"11000100",	-- 0x0B23
		"11000010",	-- 0x0B24
		"11001101",	-- 0x0B25
		"00101010",	-- 0x0B26
		"11000001",	-- 0x0B27
		"11001011",	-- 0x0B28
		"01000110",	-- 0x0B29
		"00101000",	-- 0x0B2A
		"00000100",	-- 0x0B2B
		"00011011",	-- 0x0B2C
		"11001101",	-- 0x0B2D
		"00101010",	-- 0x0B2E
		"11000001",	-- 0x0B2F
		"00011011",	-- 0x0B30
		"11001101",	-- 0x0B31
		"01000100",	-- 0x0B32
		"11000011",	-- 0x0B33
		"11001011",	-- 0x0B34
		"01111110",	-- 0x0B35
		"11000100",	-- 0x0B36
		"01001000",	-- 0x0B37
		"11000011",	-- 0x0B38
		"00100011",	-- 0x0B39
		"00011000",	-- 0x0B3A
		"11100001",	-- 0x0B3B
		"01111110",	-- 0x0B3C
		"11001101",	-- 0x0B3D
		"00110111",	-- 0x0B3E
		"11000001",	-- 0x0B3F
		"00100011",	-- 0x0B40
		"00010000",	-- 0x0B41
		"11111001",	-- 0x0B42
		"11001001",	-- 0x0B43
		"00111110",	-- 0x0B44
		"00100000",	-- 0x0B45
		"00011000",	-- 0x0B46
		"00000010",	-- 0x0B47
		"00111110",	-- 0x0B48
		"00001101",	-- 0x0B49
		"11000011",	-- 0x0B4A
		"00110111",	-- 0x0B4B
		"11000001",	-- 0x0B4C
		"01010011",	-- 0x0B4D
		"01010000",	-- 0x0B4E
		"00000001",	-- 0x0B4F
		"01010000",	-- 0x0B50
		"01000011",	-- 0x0B51
		"10000001",	-- 0x0B52
		"01000001",	-- 0x0B53
		"00110001",	-- 0x0B54
		"00000000",	-- 0x0B55
		"01000110",	-- 0x0B56
		"00110001",	-- 0x0B57
		"00000000",	-- 0x0B58
		"01000010",	-- 0x0B59
		"00110001",	-- 0x0B5A
		"00000000",	-- 0x0B5B
		"01000011",	-- 0x0B5C
		"00110001",	-- 0x0B5D
		"00000000",	-- 0x0B5E
		"01000100",	-- 0x0B5F
		"00110001",	-- 0x0B60
		"00000000",	-- 0x0B61
		"01000101",	-- 0x0B62
		"00110001",	-- 0x0B63
		"00000000",	-- 0x0B64
		"01001000",	-- 0x0B65
		"00110001",	-- 0x0B66
		"00000000",	-- 0x0B67
		"01001100",	-- 0x0B68
		"00110001",	-- 0x0B69
		"10000000",	-- 0x0B6A
		"01000001",	-- 0x0B6B
		"00110010",	-- 0x0B6C
		"00000000",	-- 0x0B6D
		"01000110",	-- 0x0B6E
		"00110010",	-- 0x0B6F
		"00000000",	-- 0x0B70
		"01000010",	-- 0x0B71
		"00110010",	-- 0x0B72
		"00000000",	-- 0x0B73
		"01000011",	-- 0x0B74
		"00110010",	-- 0x0B75
		"00000000",	-- 0x0B76
		"01000100",	-- 0x0B77
		"00110010",	-- 0x0B78
		"00000000",	-- 0x0B79
		"01000101",	-- 0x0B7A
		"00110010",	-- 0x0B7B
		"00000000",	-- 0x0B7C
		"01001000",	-- 0x0B7D
		"00110010",	-- 0x0B7E
		"00000000",	-- 0x0B7F
		"01001100",	-- 0x0B80
		"00110010",	-- 0x0B81
		"10000000",	-- 0x0B82
		"01001001",	-- 0x0B83
		"01011000",	-- 0x0B84
		"00000001",	-- 0x0B85
		"01001001",	-- 0x0B86
		"01011001",	-- 0x0B87
		"00000001",	-- 0x0B88
		"01001001",	-- 0x0B89
		"01010010",	-- 0x0B8A
		"00000000",	-- 0x0B8B
		"00000000",	-- 0x0B8C
		"11001101",	-- 0x0B8D
		"10010101",	-- 0x0B8E
		"11000001",	-- 0x0B8F
		"11110101",	-- 0x0B90
		"01111010",	-- 0x0B91
		"11111110",	-- 0x0B92
		"00001101",	-- 0x0B93
		"11000010",	-- 0x0B94
		"11111001",	-- 0x0B95
		"11000000",	-- 0x0B96
		"11110001",	-- 0x0B97
		"00110000",	-- 0x0B98
		"00000100",	-- 0x0B99
		"11101101",	-- 0x0B9A
		"01000011",	-- 0x0B9B
		"01010110",	-- 0x0B9C
		"11111100",	-- 0x0B9D
		"11110011",	-- 0x0B9E
		"00110001",	-- 0x0B9F
		"01000000",	-- 0x0BA0
		"11111100",	-- 0x0BA1
		"00111010",	-- 0x0BA2
		"01011011",	-- 0x0BA3
		"11111100",	-- 0x0BA4
		"11001011",	-- 0x0BA5
		"10000111",	-- 0x0BA6
		"00110010",	-- 0x0BA7
		"01011011",	-- 0x0BA8
		"11111100",	-- 0x0BA9
		"10101111",	-- 0x0BAA
		"11110001",	-- 0x0BAB
		"11101101",	-- 0x0BAC
		"01000111",	-- 0x0BAD
		"11111101",	-- 0x0BAE
		"11100001",	-- 0x0BAF
		"11011101",	-- 0x0BB0
		"11100001",	-- 0x0BB1
		"11100001",	-- 0x0BB2
		"11010001",	-- 0x0BB3
		"11000001",	-- 0x0BB4
		"11110001",	-- 0x0BB5
		"11011001",	-- 0x0BB6
		"00001000",	-- 0x0BB7
		"11100001",	-- 0x0BB8
		"11010001",	-- 0x0BB9
		"11000001",	-- 0x0BBA
		"11000011",	-- 0x0BBB
		"11110101",	-- 0x0BBC
		"11111100",	-- 0x0BBD
		"11110001",	-- 0x0BBE
		"11101101",	-- 0x0BBF
		"01111011",	-- 0x0BC0
		"01011000",	-- 0x0BC1
		"11111100",	-- 0x0BC2
		"00101010",	-- 0x0BC3
		"01010110",	-- 0x0BC4
		"11111100",	-- 0x0BC5
		"11100101",	-- 0x0BC6
		"00101010",	-- 0x0BC7
		"01001110",	-- 0x0BC8
		"11111100",	-- 0x0BC9
		"11111011",	-- 0x0BCA
		"11001001",	-- 0x0BCB
		"11001101",	-- 0x0BCC
		"10010101",	-- 0x0BCD
		"11000001",	-- 0x0BCE
		"11101101",	-- 0x0BCF
		"01111000",	-- 0x0BD0
		"11001101",	-- 0x0BD1
		"00101011",	-- 0x0BD2
		"11000001",	-- 0x0BD3
		"11000011",	-- 0x0BD4
		"01100001",	-- 0x0BD5
		"11000010",	-- 0x0BD6
		"11001101",	-- 0x0BD7
		"01100111",	-- 0x0BD8
		"11000010",	-- 0x0BD9
		"01001101",	-- 0x0BDA
		"11101101",	-- 0x0BDB
		"01011001",	-- 0x0BDC
		"11000011",	-- 0x0BDD
		"01100001",	-- 0x0BDE
		"11000010",	-- 0x0BDF
		"11111110",	-- 0x0BE0
		"01000001",	-- 0x0BE1
		"11011000",	-- 0x0BE2
		"11111110",	-- 0x0BE3
		"01011011",	-- 0x0BE4
		"11011000",	-- 0x0BE5
		"11111110",	-- 0x0BE6
		"01100001",	-- 0x0BE7
		"11011000",	-- 0x0BE8
		"11111110",	-- 0x0BE9
		"01111011",	-- 0x0BEA
		"11010000",	-- 0x0BEB
		"11001011",	-- 0x0BEC
		"10101111",	-- 0x0BED
		"11001001",	-- 0x0BEE
		"00100001",	-- 0x0BEF
		"00101010",	-- 0x0BF0
		"11000100",	-- 0x0BF1
		"00100010",	-- 0x0BF2
		"00000000",	-- 0x0BF3
		"11111101",	-- 0x0BF4
		"11001101",	-- 0x0BF5
		"11010001",	-- 0x0BF6
		"11000101",	-- 0x0BF7
		"10101111",	-- 0x0BF8
		"00110010",	-- 0x0BF9
		"01011101",	-- 0x0BFA
		"11111100",	-- 0x0BFB
		"00100001",	-- 0x0BFC
		"00001100",	-- 0x0BFD
		"11000100",	-- 0x0BFE
		"00001110",	-- 0x0BFF
		"11100111",	-- 0x0C00
		"00000110",	-- 0x0C01
		"00001100",	-- 0x0C02
		"11101101",	-- 0x0C03
		"10110011",	-- 0x0C04
		"00000110",	-- 0x0C05
		"00000010",	-- 0x0C06
		"00001110",	-- 0x0C07
		"11110100",	-- 0x0C08
		"11101101",	-- 0x0C09
		"10110011",	-- 0x0C0A
		"11001001",	-- 0x0C0B
		"00000000",	-- 0x0C0C
		"00011000",	-- 0x0C0D
		"00000001",	-- 0x0C0E
		"00011000",	-- 0x0C0F
		"00000010",	-- 0x0C10
		"00000000",	-- 0x0C11
		"00000011",	-- 0x0C12
		"11000001",	-- 0x0C13
		"00000100",	-- 0x0C14
		"01000100",	-- 0x0C15
		"00000101",	-- 0x0C16
		"01101000",	-- 0x0C17
		"01000111",	-- 0x0C18
		"00001101",	-- 0x0C19
		"11000011",	-- 0x0C1A
		"11111100",	-- 0x0C1B
		"11111100",	-- 0x0C1C
		"00111010",	-- 0x0C1D
		"01011010",	-- 0x0C1E
		"11111100",	-- 0x0C1F
		"10110111",	-- 0x0C20
		"00101000",	-- 0x0C21
		"11110111",	-- 0x0C22
		"11110101",	-- 0x0C23
		"10101111",	-- 0x0C24
		"00110010",	-- 0x0C25
		"01011010",	-- 0x0C26
		"11111100",	-- 0x0C27
		"11110001",	-- 0x0C28
		"11001001",	-- 0x0C29
		"11110101",	-- 0x0C2A
		"11011011",	-- 0x0C2B
		"11100101",	-- 0x0C2C
		"00110010",	-- 0x0C2D
		"01011010",	-- 0x0C2E
		"11111100",	-- 0x0C2F
		"11110001",	-- 0x0C30
		"11111011",	-- 0x0C31
		"11101101",	-- 0x0C32
		"01001101",	-- 0x0C33
		"01001111",	-- 0x0C34
		"11110101",	-- 0x0C35
		"00111010",	-- 0x0C36
		"01011011",	-- 0x0C37
		"11111100",	-- 0x0C38
		"11001011",	-- 0x0C39
		"01001111",	-- 0x0C3A
		"00100000",	-- 0x0C3B
		"11111001",	-- 0x0C3C
		"11110001",	-- 0x0C3D
		"11000011",	-- 0x0C3E
		"11111001",	-- 0x0C3F
		"11111100",	-- 0x0C40
		"00100001",	-- 0x0C41
		"01011110",	-- 0x0C42
		"11111100",	-- 0x0C43
		"00010110",	-- 0x0C44
		"00000000",	-- 0x0C45
		"01000110",	-- 0x0C46
		"00100011",	-- 0x0C47
		"00001110",	-- 0x0C48
		"11111001",	-- 0x0C49
		"11001101",	-- 0x0C4A
		"01101010",	-- 0x0C4B
		"11000100",	-- 0x0C4C
		"00100000",	-- 0x0C4D
		"00010100",	-- 0x0C4E
		"11101101",	-- 0x0C4F
		"10100011",	-- 0x0C50
		"00100000",	-- 0x0C51
		"11110111",	-- 0x0C52
		"00100001",	-- 0x0C53
		"01101001",	-- 0x0C54
		"11111100",	-- 0x0C55
		"11001101",	-- 0x0C56
		"01101010",	-- 0x0C57
		"11000100",	-- 0x0C58
		"01111010",	-- 0x0C59
		"00110010",	-- 0x0C5A
		"01101000",	-- 0x0C5B
		"11111100",	-- 0x0C5C
		"11001000",	-- 0x0C5D
		"00010100",	-- 0x0C5E
		"11101101",	-- 0x0C5F
		"10100010",	-- 0x0C60
		"00011000",	-- 0x0C61
		"11110011",	-- 0x0C62
		"10101111",	-- 0x0C63
		"01010111",	-- 0x0C64
		"11001101",	-- 0x0C65
		"01010011",	-- 0x0C66
		"11000100",	-- 0x0C67
		"00110111",	-- 0x0C68
		"11001001",	-- 0x0C69
		"11011011",	-- 0x0C6A
		"11111000",	-- 0x0C6B
		"11001011",	-- 0x0C6C
		"01111111",	-- 0x0C6D
		"00101000",	-- 0x0C6E
		"11111010",	-- 0x0C6F
		"10100111",	-- 0x0C70
		"11001011",	-- 0x0C71
		"01110111",	-- 0x0C72
		"11001001",	-- 0x0C73
		"00100001",	-- 0x0C74
		"11011100",	-- 0x0C75
		"11111100",	-- 0x0C76
		"00100010",	-- 0x0C77
		"00100000",	-- 0x0C78
		"11111101",	-- 0x0C79
		"11011011",	-- 0x0C7A
		"11101100",	-- 0x0C7B
		"11110110",	-- 0x0C7C
		"00000001",	-- 0x0C7D
		"11010011",	-- 0x0C7E
		"11101100",	-- 0x0C7F
		"00000001",	-- 0x0C80
		"00000000",	-- 0x0C81
		"00010000",	-- 0x0C82
		"11000101",	-- 0x0C83
		"00100001",	-- 0x0C84
		"11001000",	-- 0x0C85
		"11000100",	-- 0x0C86
		"00010001",	-- 0x0C87
		"01011110",	-- 0x0C88
		"11111100",	-- 0x0C89
		"00000001",	-- 0x0C8A
		"00000011",	-- 0x0C8B
		"00000000",	-- 0x0C8C
		"11101101",	-- 0x0C8D
		"10110000",	-- 0x0C8E
		"11001101",	-- 0x0C8F
		"01000001",	-- 0x0C90
		"11000100",	-- 0x0C91
		"00111010",	-- 0x0C92
		"01101001",	-- 0x0C93
		"11111100",	-- 0x0C94
		"11000001",	-- 0x0C95
		"11001011",	-- 0x0C96
		"01101111",	-- 0x0C97
		"11000010",	-- 0x0C98
		"10100011",	-- 0x0C99
		"11000100",	-- 0x0C9A
		"00001011",	-- 0x0C9B
		"01111000",	-- 0x0C9C
		"10110001",	-- 0x0C9D
		"11001010",	-- 0x0C9E
		"10100011",	-- 0x0C9F
		"11000101",	-- 0x0CA0
		"00011000",	-- 0x0CA1
		"11100000",	-- 0x0CA2
		"00100001",	-- 0x0CA3
		"11001011",	-- 0x0CA4
		"11000100",	-- 0x0CA5
		"00010001",	-- 0x0CA6
		"01011110",	-- 0x0CA7
		"11111100",	-- 0x0CA8
		"00000001",	-- 0x0CA9
		"00000100",	-- 0x0CAA
		"00000000",	-- 0x0CAB
		"11101101",	-- 0x0CAC
		"10110000",	-- 0x0CAD
		"11001101",	-- 0x0CAE
		"01000001",	-- 0x0CAF
		"11000100",	-- 0x0CB0
		"00100001",	-- 0x0CB1
		"11001111",	-- 0x0CB2
		"11000100",	-- 0x0CB3
		"00010001",	-- 0x0CB4
		"01011110",	-- 0x0CB5
		"11111100",	-- 0x0CB6
		"00000001",	-- 0x0CB7
		"00000011",	-- 0x0CB8
		"00000000",	-- 0x0CB9
		"11101101",	-- 0x0CBA
		"10110000",	-- 0x0CBB
		"11001101",	-- 0x0CBC
		"00001010",	-- 0x0CBD
		"11000101",	-- 0x0CBE
		"00000110",	-- 0x0CBF
		"00000110",	-- 0x0CC0
		"00111110",	-- 0x0CC1
		"11000011",	-- 0x0CC2
		"11010011",	-- 0x0CC3
		"11111111",	-- 0x0CC4
		"00010000",	-- 0x0CC5
		"11111100",	-- 0x0CC6
		"11001001",	-- 0x0CC7
		"00000010",	-- 0x0CC8
		"00000100",	-- 0x0CC9
		"00000000",	-- 0x0CCA
		"00000011",	-- 0x0CCB
		"00000011",	-- 0x0CCC
		"11110011",	-- 0x0CCD
		"11111110",	-- 0x0CCE
		"00000010",	-- 0x0CCF
		"00000111",	-- 0x0CD0
		"00000000",	-- 0x0CD1
		"01111001",	-- 0x0CD2
		"10000000",	-- 0x0CD3
		"10011111",	-- 0x0CD4
		"11111111",	-- 0x0CD5
		"00010011",	-- 0x0CD6
		"01010100",	-- 0x0CD7
		"01111100",	-- 0x0CD8
		"01101000",	-- 0x0CD9
		"10111100",	-- 0x0CDA
		"11010101",	-- 0x0CDB
		"11111101",	-- 0x0CDC
		"00010010",	-- 0x0CDD
		"00100000",	-- 0x0CDE
		"10001010",	-- 0x0CDF
		"11001111",	-- 0x0CE0
		"11100000",	-- 0x0CE1
		"00001001",	-- 0x0CE2
		"01000110",	-- 0x0CE3
		"00000000",	-- 0x0CE4
		"00000000",	-- 0x0CE5
		"00000000",	-- 0x0CE6
		"00000001",	-- 0x0CE7
		"00000011",	-- 0x0CE8
		"00000101",	-- 0x0CE9
		"00100101",	-- 0x0CEA
		"11111111",	-- 0x0CEB
		"00000011",	-- 0x0CEC
		"00001111",	-- 0x0CED
		"00000000",	-- 0x0CEE
		"00000001",	-- 0x0CEF
		"01111001",	-- 0x0CF0
		"10000000",	-- 0x0CF1
		"10110011",	-- 0x0CF2
		"01111111",	-- 0x0CF3
		"00001100",	-- 0x0CF4
		"01010100",	-- 0x0CF5
		"01111100",	-- 0x0CF6
		"01101000",	-- 0x0CF7
		"10111100",	-- 0x0CF8
		"11010101",	-- 0x0CF9
		"11111101",	-- 0x0CFA
		"00010010",	-- 0x0CFB
		"00100000",	-- 0x0CFC
		"10001010",	-- 0x0CFD
		"11001111",	-- 0x0CFE
		"11100000",	-- 0x0CFF
		"00001001",	-- 0x0D00
		"01000110",	-- 0x0D01
		"00000000",	-- 0x0D02
		"00000001",	-- 0x0D03
		"00000000",	-- 0x0D04
		"00000001",	-- 0x0D05
		"00000011",	-- 0x0D06
		"00000101",	-- 0x0D07
		"00100101",	-- 0x0D08
		"11111111",	-- 0x0D09
		"11001101",	-- 0x0D0A
		"01000001",	-- 0x0D0B
		"11000100",	-- 0x0D0C
		"11011010",	-- 0x0D0D
		"10100011",	-- 0x0D0E
		"11000101",	-- 0x0D0F
		"00111010",	-- 0x0D10
		"01101000",	-- 0x0D11
		"11111100",	-- 0x0D12
		"10110111",	-- 0x0D13
		"11000010",	-- 0x0D14
		"10100011",	-- 0x0D15
		"11000101",	-- 0x0D16
		"00111100",	-- 0x0D17
		"00110010",	-- 0x0D18
		"01011110",	-- 0x0D19
		"11111100",	-- 0x0D1A
		"00111110",	-- 0x0D1B
		"00001000",	-- 0x0D1C
		"00110010",	-- 0x0D1D
		"01011111",	-- 0x0D1E
		"11111100",	-- 0x0D1F
		"11001101",	-- 0x0D20
		"01000001",	-- 0x0D21
		"11000100",	-- 0x0D22
		"11011010",	-- 0x0D23
		"10100011",	-- 0x0D24
		"11000101",	-- 0x0D25
		"00111010",	-- 0x0D26
		"01101001",	-- 0x0D27
		"11111100",	-- 0x0D28
		"11111110",	-- 0x0D29
		"10000000",	-- 0x0D2A
		"00101000",	-- 0x0D2B
		"11110011",	-- 0x0D2C
		"11100110",	-- 0x0D2D
		"11100000",	-- 0x0D2E
		"11111110",	-- 0x0D2F
		"00100000",	-- 0x0D30
		"00001111",	-- 0x0D31
		"11001000",	-- 0x0D32
		"11000011",	-- 0x0D33
		"10100011",	-- 0x0D34
		"11000101",	-- 0x0D35
		"00000110",	-- 0x0D36
		"00001010",	-- 0x0D37
		"11000101",	-- 0x0D38
		"11001101",	-- 0x0D39
		"01110100",	-- 0x0D3A
		"11000100",	-- 0x0D3B
		"00100001",	-- 0x0D3C
		"11010010",	-- 0x0D3D
		"11000100",	-- 0x0D3E
		"00001110",	-- 0x0D3F
		"11111111",	-- 0x0D40
		"00000110",	-- 0x0D41
		"00010000",	-- 0x0D42
		"11101101",	-- 0x0D43
		"10110011",	-- 0x0D44
		"00100001",	-- 0x0D45
		"11100010",	-- 0x0D46
		"11000100",	-- 0x0D47
		"00010001",	-- 0x0D48
		"01011110",	-- 0x0D49
		"11111100",	-- 0x0D4A
		"00000001",	-- 0x0D4B
		"00001010",	-- 0x0D4C
		"00000000",	-- 0x0D4D
		"11101101",	-- 0x0D4E
		"10110000",	-- 0x0D4F
		"11001101",	-- 0x0D50
		"01000001",	-- 0x0D51
		"11000100",	-- 0x0D52
		"00111010",	-- 0x0D53
		"01101000",	-- 0x0D54
		"11111100",	-- 0x0D55
		"11111110",	-- 0x0D56
		"00000111",	-- 0x0D57
		"00100000",	-- 0x0D58
		"01001010",	-- 0x0D59
		"00111010",	-- 0x0D5A
		"01101001",	-- 0x0D5B
		"11111100",	-- 0x0D5C
		"11100110",	-- 0x0D5D
		"11000000",	-- 0x0D5E
		"00100000",	-- 0x0D5F
		"01000011",	-- 0x0D60
		"00100001",	-- 0x0D61
		"11101100",	-- 0x0D62
		"11000100",	-- 0x0D63
		"00010001",	-- 0x0D64
		"01011110",	-- 0x0D65
		"11111100",	-- 0x0D66
		"00000001",	-- 0x0D67
		"00000100",	-- 0x0D68
		"00000000",	-- 0x0D69
		"11101101",	-- 0x0D6A
		"10110000",	-- 0x0D6B
		"11001101",	-- 0x0D6C
		"00001010",	-- 0x0D6D
		"11000101",	-- 0x0D6E
		"00100001",	-- 0x0D6F
		"11110000",	-- 0x0D70
		"11000100",	-- 0x0D71
		"00001110",	-- 0x0D72
		"11111111",	-- 0x0D73
		"00000110",	-- 0x0D74
		"00010000",	-- 0x0D75
		"11101101",	-- 0x0D76
		"10110011",	-- 0x0D77
		"00100001",	-- 0x0D78
		"00000000",	-- 0x0D79
		"11000101",	-- 0x0D7A
		"00010001",	-- 0x0D7B
		"01011110",	-- 0x0D7C
		"11111100",	-- 0x0D7D
		"00000001",	-- 0x0D7E
		"00001010",	-- 0x0D7F
		"00000000",	-- 0x0D80
		"11101101",	-- 0x0D81
		"10110000",	-- 0x0D82
		"11001101",	-- 0x0D83
		"01000001",	-- 0x0D84
		"11000100",	-- 0x0D85
		"00111010",	-- 0x0D86
		"01101000",	-- 0x0D87
		"11111100",	-- 0x0D88
		"11111110",	-- 0x0D89
		"00000111",	-- 0x0D8A
		"00100000",	-- 0x0D8B
		"00010111",	-- 0x0D8C
		"00111010",	-- 0x0D8D
		"01101001",	-- 0x0D8E
		"11111100",	-- 0x0D8F
		"11100110",	-- 0x0D90
		"11000000",	-- 0x0D91
		"00100000",	-- 0x0D92
		"00010000",	-- 0x0D93
		"11001101",	-- 0x0D94
		"01001000",	-- 0x0D95
		"11000011",	-- 0x0D96
		"00111010",	-- 0x0D97
		"01011011",	-- 0x0D98
		"11111100",	-- 0x0D99
		"11001011",	-- 0x0D9A
		"10000111",	-- 0x0D9B
		"00110010",	-- 0x0D9C
		"01011011",	-- 0x0D9D
		"11111100",	-- 0x0D9E
		"11000001",	-- 0x0D9F
		"11000011",	-- 0x0DA0
		"10000000",	-- 0x0DA1
		"10011111",	-- 0x0DA2
		"11100001",	-- 0x0DA3
		"11000001",	-- 0x0DA4
		"00010000",	-- 0x0DA5
		"10010001",	-- 0x0DA6
		"11011011",	-- 0x0DA7
		"11101100",	-- 0x0DA8
		"11101110",	-- 0x0DA9
		"00000001",	-- 0x0DAA
		"11010011",	-- 0x0DAB
		"11101100",	-- 0x0DAC
		"11000011",	-- 0x0DAD
		"11111001",	-- 0x0DAE
		"11000000",	-- 0x0DAF
		"11110101",	-- 0x0DB0
		"00111110",	-- 0x0DB1
		"10100011",	-- 0x0DB2
		"11010011",	-- 0x0DB3
		"11111111",	-- 0x0DB4
		"11110001",	-- 0x0DB5
		"11111011",	-- 0x0DB6
		"11101101",	-- 0x0DB7
		"01001101",	-- 0x0DB8
		"00111010",	-- 0x0DB9
		"01011010",	-- 0x0DBA
		"11111100",	-- 0x0DBB
		"10110111",	-- 0x0DBC
		"00101000",	-- 0x0DBD
		"00000010",	-- 0x0DBE
		"00111110",	-- 0x0DBF
		"11111111",	-- 0x0DC0
		"11111110",	-- 0x0DC1
		"11111111",	-- 0x0DC2
		"11001001",	-- 0x0DC3
		"00000000",	-- 0x0DC4
		"11110101",	-- 0x0DC5
		"11000101",	-- 0x0DC6
		"11010101",	-- 0x0DC7
		"11100101",	-- 0x0DC8
		"11001101",	-- 0x0DC9
		"11000110",	-- 0x0DCA
		"11000111",	-- 0x0DCB
		"11100001",	-- 0x0DCC
		"11010001",	-- 0x0DCD
		"11000001",	-- 0x0DCE
		"11110001",	-- 0x0DCF
		"11001001",	-- 0x0DD0
		"11110101",	-- 0x0DD1
		"11000101",	-- 0x0DD2
		"11010101",	-- 0x0DD3
		"11100101",	-- 0x0DD4
		"11001101",	-- 0x0DD5
		"11111011",	-- 0x0DD6
		"11000101",	-- 0x0DD7
		"11001101",	-- 0x0DD8
		"01010111",	-- 0x0DD9
		"11001000",	-- 0x0DDA
		"00111110",	-- 0x0DDB
		"00011011",	-- 0x0DDC
		"00110010",	-- 0x0DDD
		"00100110",	-- 0x0DDE
		"11111100",	-- 0x0DDF
		"00011000",	-- 0x0DE0
		"11101010",	-- 0x0DE1
		"00001000",	-- 0x0DE2
		"00010110",	-- 0x0DE3
		"00101100",	-- 0x0DE4
		"10000101",	-- 0x0DE5
		"00010101",	-- 0x0DE6
		"00000101",	-- 0x0DE7
		"00000010",	-- 0x0DE8
		"00001000",	-- 0x0DE9
		"01111101",	-- 0x0DEA
		"00001000",	-- 0x0DEB
		"00010110",	-- 0x0DEC
		"00101100",	-- 0x0DED
		"10000101",	-- 0x0DEE
		"00000101",	-- 0x0DEF
		"00000001",	-- 0x0DF0
		"00101111",	-- 0x0DF1
		"00001000",	-- 0x0DF2
		"11000001",	-- 0x0DF3
		"00000110",	-- 0x0DF4
		"10000000",	-- 0x0DF5
		"00010000",	-- 0x0DF6
		"00000000",	-- 0x0DF7
		"00000000",	-- 0x0DF8
		"00000000",	-- 0x0DF9
		"00000000",	-- 0x0DFA
		"10101111",	-- 0x0DFB
		"00110010",	-- 0x0DFC
		"00001001",	-- 0x0DFD
		"11111100",	-- 0x0DFE
		"00110010",	-- 0x0DFF
		"00001001",	-- 0x0E00
		"11111100",	-- 0x0E01
		"00110010",	-- 0x0E02
		"00010101",	-- 0x0E03
		"11111100",	-- 0x0E04
		"00111100",	-- 0x0E05
		"00110010",	-- 0x0E06
		"00000000",	-- 0x0E07
		"11111100",	-- 0x0E08
		"00110010",	-- 0x0E09
		"00010110",	-- 0x0E0A
		"11111100",	-- 0x0E0B
		"00110010",	-- 0x0E0C
		"00011100",	-- 0x0E0D
		"11111100",	-- 0x0E0E
		"00110010",	-- 0x0E0F
		"00000001",	-- 0x0E10
		"11111100",	-- 0x0E11
		"00111110",	-- 0x0E12
		"00000000",	-- 0x0E13
		"11010011",	-- 0x0E14
		"01110001",	-- 0x0E15
		"00001110",	-- 0x0E16
		"01110000",	-- 0x0E17
		"00100001",	-- 0x0E18
		"11100010",	-- 0x0E19
		"11000101",	-- 0x0E1A
		"11011011",	-- 0x0E1B
		"11100111",	-- 0x0E1C
		"11001011",	-- 0x0E1D
		"01101111",	-- 0x0E1E
		"00101000",	-- 0x0E1F
		"00000011",	-- 0x0E20
		"00100001",	-- 0x0E21
		"11101011",	-- 0x0E22
		"11000101",	-- 0x0E23
		"01000110",	-- 0x0E24
		"00100011",	-- 0x0E25
		"11101101",	-- 0x0E26
		"10110011",	-- 0x0E27
		"11001101",	-- 0x0E28
		"11000100",	-- 0x0E29
		"11000110",	-- 0x0E2A
		"00111110",	-- 0x0E2B
		"01101111",	-- 0x0E2C
		"11010011",	-- 0x0E2D
		"01110001",	-- 0x0E2E
		"00100001",	-- 0x0E2F
		"11110100",	-- 0x0E30
		"11000101",	-- 0x0E31
		"01000110",	-- 0x0E32
		"00100011",	-- 0x0E33
		"00111110",	-- 0x0E34
		"01110010",	-- 0x0E35
		"11010011",	-- 0x0E36
		"01110001",	-- 0x0E37
		"11101101",	-- 0x0E38
		"10110011",	-- 0x0E39
		"00111110",	-- 0x0E3A
		"01001010",	-- 0x0E3B
		"11010011",	-- 0x0E3C
		"01110001",	-- 0x0E3D
		"00111110",	-- 0x0E3E
		"11111111",	-- 0x0E3F
		"11101101",	-- 0x0E40
		"01111001",	-- 0x0E41
		"11101101",	-- 0x0E42
		"01111001",	-- 0x0E43
		"00111110",	-- 0x0E44
		"01000111",	-- 0x0E45
		"11010011",	-- 0x0E46
		"01110001",	-- 0x0E47
		"00111110",	-- 0x0E48
		"00101110",	-- 0x0E49
		"11101101",	-- 0x0E4A
		"01111001",	-- 0x0E4B
		"00100001",	-- 0x0E4C
		"00000000",	-- 0x0E4D
		"00000000",	-- 0x0E4E
		"00100010",	-- 0x0E4F
		"00000101",	-- 0x0E50
		"11111100",	-- 0x0E51
		"11001101",	-- 0x0E52
		"10110100",	-- 0x0E53
		"11000110",	-- 0x0E54
		"00010001",	-- 0x0E55
		"00000111",	-- 0x0E56
		"00000001",	-- 0x0E57
		"00100001",	-- 0x0E58
		"01000010",	-- 0x0E59
		"00101111",	-- 0x0E5A
		"11101101",	-- 0x0E5B
		"01001011",	-- 0x0E5C
		"00000101",	-- 0x0E5D
		"11111100",	-- 0x0E5E
		"00001001",	-- 0x0E5F
		"00100010",	-- 0x0E60
		"00000010",	-- 0x0E61
		"11111100",	-- 0x0E62
		"10101111",	-- 0x0E63
		"00110010",	-- 0x0E64
		"00000100",	-- 0x0E65
		"11111100",	-- 0x0E66
		"11001101",	-- 0x0E67
		"01111111",	-- 0x0E68
		"11000111",	-- 0x0E69
		"00111110",	-- 0x0E6A
		"00110000",	-- 0x0E6B
		"11010011",	-- 0x0E6C
		"01110001",	-- 0x0E6D
		"11001101",	-- 0x0E6E
		"11000100",	-- 0x0E6F
		"11000110",	-- 0x0E70
		"00111110",	-- 0x0E71
		"01001100",	-- 0x0E72
		"11010011",	-- 0x0E73
		"01110001",	-- 0x0E74
		"00111110",	-- 0x0E75
		"00010010",	-- 0x0E76
		"11101101",	-- 0x0E77
		"01111001",	-- 0x0E78
		"11101101",	-- 0x0E79
		"01011001",	-- 0x0E7A
		"11101101",	-- 0x0E7B
		"01010001",	-- 0x0E7C
		"00100001",	-- 0x0E7D
		"11100000",	-- 0x0E7E
		"00000010",	-- 0x0E7F
		"11101101",	-- 0x0E80
		"01101001",	-- 0x0E81
		"11101101",	-- 0x0E82
		"01100001",	-- 0x0E83
		"11101101",	-- 0x0E84
		"01101001",	-- 0x0E85
		"11101101",	-- 0x0E86
		"01100001",	-- 0x0E87
		"11001101",	-- 0x0E88
		"11000100",	-- 0x0E89
		"11000110",	-- 0x0E8A
		"00111110",	-- 0x0E8B
		"01000110",	-- 0x0E8C
		"11010011",	-- 0x0E8D
		"01110001",	-- 0x0E8E
		"10101111",	-- 0x0E8F
		"11101101",	-- 0x0E90
		"01111001",	-- 0x0E91
		"00111110",	-- 0x0E92
		"01111000",	-- 0x0E93
		"11010011",	-- 0x0E94
		"01110001",	-- 0x0E95
		"00000110",	-- 0x0E96
		"00001000",	-- 0x0E97
		"00111110",	-- 0x0E98
		"00000000",	-- 0x0E99
		"11101101",	-- 0x0E9A
		"01111001",	-- 0x0E9B
		"00010000",	-- 0x0E9C
		"11111100",	-- 0x0E9D
		"00100001",	-- 0x0E9E
		"01101000",	-- 0x0E9F
		"00001101",	-- 0x0EA0
		"00001110",	-- 0x0EA1
		"01110001",	-- 0x0EA2
		"11101101",	-- 0x0EA3
		"01101001",	-- 0x0EA4
		"11101101",	-- 0x0EA5
		"01100001",	-- 0x0EA6
		"00111110",	-- 0x0EA7
		"00000001",	-- 0x0EA8
		"00110010",	-- 0x0EA9
		"00000000",	-- 0x0EAA
		"11111100",	-- 0x0EAB
		"00111110",	-- 0x0EAC
		"00000001",	-- 0x0EAD
		"00110010",	-- 0x0EAE
		"00000001",	-- 0x0EAF
		"11111100",	-- 0x0EB0
		"11000011",	-- 0x0EB1
		"00101101",	-- 0x0EB2
		"11000111",	-- 0x0EB3
		"11001101",	-- 0x0EB4
		"11000100",	-- 0x0EB5
		"11000110",	-- 0x0EB6
		"00111110",	-- 0x0EB7
		"01110000",	-- 0x0EB8
		"00100001",	-- 0x0EB9
		"00000101",	-- 0x0EBA
		"11111100",	-- 0x0EBB
		"11010011",	-- 0x0EBC
		"01110001",	-- 0x0EBD
		"00000001",	-- 0x0EBE
		"01110000",	-- 0x0EBF
		"00000010",	-- 0x0EC0
		"11101101",	-- 0x0EC1
		"10110011",	-- 0x0EC2
		"11001001",	-- 0x0EC3
		"11011011",	-- 0x0EC4
		"01110000",	-- 0x0EC5
		"11001011",	-- 0x0EC6
		"01010111",	-- 0x0EC7
		"11000000",	-- 0x0EC8
		"00011000",	-- 0x0EC9
		"11111001",	-- 0x0ECA
		"11011011",	-- 0x0ECB
		"01110000",	-- 0x0ECC
		"11001011",	-- 0x0ECD
		"01001111",	-- 0x0ECE
		"11001000",	-- 0x0ECF
		"00011000",	-- 0x0ED0
		"11111001",	-- 0x0ED1
		"11011011",	-- 0x0ED2
		"01110000",	-- 0x0ED3
		"11001011",	-- 0x0ED4
		"01000111",	-- 0x0ED5
		"11001001",	-- 0x0ED6
		"00010110",	-- 0x0ED7
		"00000001",	-- 0x0ED8
		"00011110",	-- 0x0ED9
		"00001001",	-- 0x0EDA
		"11001101",	-- 0x0EDB
		"11000100",	-- 0x0EDC
		"11000110",	-- 0x0EDD
		"00111110",	-- 0x0EDE
		"01000110",	-- 0x0EDF
		"11010011",	-- 0x0EE0
		"01110001",	-- 0x0EE1
		"00111110",	-- 0x0EE2
		"00000001",	-- 0x0EE3
		"00111101",	-- 0x0EE4
		"11010011",	-- 0x0EE5
		"01110000",	-- 0x0EE6
		"00111110",	-- 0x0EE7
		"01001100",	-- 0x0EE8
		"11010011",	-- 0x0EE9
		"01110001",	-- 0x0EEA
		"00001110",	-- 0x0EEB
		"01110000",	-- 0x0EEC
		"00111110",	-- 0x0EED
		"00010010",	-- 0x0EEE
		"11101101",	-- 0x0EEF
		"01111001",	-- 0x0EF0
		"10101111",	-- 0x0EF1
		"11101101",	-- 0x0EF2
		"01010001",	-- 0x0EF3
		"11101101",	-- 0x0EF4
		"01111001",	-- 0x0EF5
		"11101101",	-- 0x0EF6
		"01011001",	-- 0x0EF7
		"11101101",	-- 0x0EF8
		"01111001",	-- 0x0EF9
		"11101101",	-- 0x0EFA
		"01011001",	-- 0x0EFB
		"11101101",	-- 0x0EFC
		"01111001",	-- 0x0EFD
		"11001101",	-- 0x0EFE
		"11000100",	-- 0x0EFF
		"11000110",	-- 0x0F00
		"00111110",	-- 0x0F01
		"01111000",	-- 0x0F02
		"11010011",	-- 0x0F03
		"01110001",	-- 0x0F04
		"00000110",	-- 0x0F05
		"00001000",	-- 0x0F06
		"00111110",	-- 0x0F07
		"11111111",	-- 0x0F08
		"11101101",	-- 0x0F09
		"01111001",	-- 0x0F0A
		"00010000",	-- 0x0F0B
		"11111100",	-- 0x0F0C
		"11001101",	-- 0x0F0D
		"11001011",	-- 0x0F0E
		"11000110",	-- 0x0F0F
		"00111110",	-- 0x0F10
		"00110001",	-- 0x0F11
		"11010011",	-- 0x0F12
		"01110001",	-- 0x0F13
		"00111110",	-- 0x0F14
		"01101000",	-- 0x0F15
		"11010011",	-- 0x0F16
		"01110001",	-- 0x0F17
		"11001001",	-- 0x0F18
		"00100001",	-- 0x0F19
		"00000000",	-- 0x0F1A
		"00000000",	-- 0x0F1B
		"00111110",	-- 0x0F1C
		"00010001",	-- 0x0F1D
		"11001011",	-- 0x0F1E
		"00011000",	-- 0x0F1F
		"11001011",	-- 0x0F20
		"00011001",	-- 0x0F21
		"00111101",	-- 0x0F22
		"11001000",	-- 0x0F23
		"00110000",	-- 0x0F24
		"00000001",	-- 0x0F25
		"00011001",	-- 0x0F26
		"11001011",	-- 0x0F27
		"00011100",	-- 0x0F28
		"11001011",	-- 0x0F29
		"00011101",	-- 0x0F2A
		"00011000",	-- 0x0F2B
		"11110001",	-- 0x0F2C
		"00010001",	-- 0x0F2D
		"00001011",	-- 0x0F2E
		"00000000",	-- 0x0F2F
		"00000001",	-- 0x0F30
		"00101110",	-- 0x0F31
		"00000000",	-- 0x0F32
		"11001101",	-- 0x0F33
		"00011001",	-- 0x0F34
		"11000111",	-- 0x0F35
		"11101101",	-- 0x0F36
		"01011011",	-- 0x0F37
		"00000000",	-- 0x0F38
		"11111100",	-- 0x0F39
		"00010110",	-- 0x0F3A
		"00000000",	-- 0x0F3B
		"11001101",	-- 0x0F3C
		"00011001",	-- 0x0F3D
		"11000111",	-- 0x0F3E
		"01100000",	-- 0x0F3F
		"01101001",	-- 0x0F40
		"00000001",	-- 0x0F41
		"00101110",	-- 0x0F42
		"00000000",	-- 0x0F43
		"10100111",	-- 0x0F44
		"11101101",	-- 0x0F45
		"01000010",	-- 0x0F46
		"11101101",	-- 0x0F47
		"01001011",	-- 0x0F48
		"00000101",	-- 0x0F49
		"11111100",	-- 0x0F4A
		"00001001",	-- 0x0F4B
		"00100010",	-- 0x0F4C
		"00000111",	-- 0x0F4D
		"11111100",	-- 0x0F4E
		"10101111",	-- 0x0F4F
		"00011110",	-- 0x0F50
		"00001001",	-- 0x0F51
		"01010111",	-- 0x0F52
		"11101101",	-- 0x0F53
		"01001011",	-- 0x0F54
		"00000001",	-- 0x0F55
		"11111100",	-- 0x0F56
		"01000111",	-- 0x0F57
		"11001101",	-- 0x0F58
		"00011001",	-- 0x0F59
		"11000111",	-- 0x0F5A
		"01100000",	-- 0x0F5B
		"01101001",	-- 0x0F5C
		"10101111",	-- 0x0F5D
		"10101111",	-- 0x0F5E
		"11101101",	-- 0x0F5F
		"01010010",	-- 0x0F60
		"00100010",	-- 0x0F61
		"00011010",	-- 0x0F62
		"11111100",	-- 0x0F63
		"00000110",	-- 0x0F64
		"00000100",	-- 0x0F65
		"11001011",	-- 0x0F66
		"00111100",	-- 0x0F67
		"11001011",	-- 0x0F68
		"00011101",	-- 0x0F69
		"11001011",	-- 0x0F6A
		"00011111",	-- 0x0F6B
		"00010000",	-- 0x0F6C
		"11111000",	-- 0x0F6D
		"00110010",	-- 0x0F6E
		"00000100",	-- 0x0F6F
		"11111100",	-- 0x0F70
		"00110010",	-- 0x0F71
		"00011001",	-- 0x0F72
		"11111100",	-- 0x0F73
		"11101101",	-- 0x0F74
		"01011011",	-- 0x0F75
		"00000111",	-- 0x0F76
		"11111100",	-- 0x0F77
		"00011001",	-- 0x0F78
		"00100010",	-- 0x0F79
		"00000010",	-- 0x0F7A
		"11111100",	-- 0x0F7B
		"00100010",	-- 0x0F7C
		"00010111",	-- 0x0F7D
		"11111100",	-- 0x0F7E
		"11001101",	-- 0x0F7F
		"11000100",	-- 0x0F80
		"11000110",	-- 0x0F81
		"00111110",	-- 0x0F82
		"01001001",	-- 0x0F83
		"00100001",	-- 0x0F84
		"00000010",	-- 0x0F85
		"11111100",	-- 0x0F86
		"11001101",	-- 0x0F87
		"10111100",	-- 0x0F88
		"11000110",	-- 0x0F89
		"00111010",	-- 0x0F8A
		"00000100",	-- 0x0F8B
		"11111100",	-- 0x0F8C
		"11100110",	-- 0x0F8D
		"11110000",	-- 0x0F8E
		"11101101",	-- 0x0F8F
		"01111001",	-- 0x0F90
		"11001001",	-- 0x0F91
		"01111001",	-- 0x0F92
		"00100001",	-- 0x0F93
		"10111010",	-- 0x0F94
		"11000111",	-- 0x0F95
		"00000001",	-- 0x0F96
		"00000100",	-- 0x0F97
		"00000000",	-- 0x0F98
		"11101101",	-- 0x0F99
		"10110001",	-- 0x0F9A
		"11000000",	-- 0x0F9B
		"11000101",	-- 0x0F9C
		"11001101",	-- 0x0F9D
		"01101000",	-- 0x0F9E
		"11001000",	-- 0x0F9F
		"11001101",	-- 0x0FA0
		"01111111",	-- 0x0FA1
		"11000111",	-- 0x0FA2
		"11000001",	-- 0x0FA3
		"00100001",	-- 0x0FA4
		"10111110",	-- 0x0FA5
		"11000111",	-- 0x0FA6
		"11001101",	-- 0x0FA7
		"10110011",	-- 0x0FA8
		"11000111",	-- 0x0FA9
		"00101010",	-- 0x0FAA
		"00011010",	-- 0x0FAB
		"11111100",	-- 0x0FAC
		"11001101",	-- 0x0FAD
		"01100001",	-- 0x0FAE
		"11000111",	-- 0x0FAF
		"11000011",	-- 0x0FB0
		"01010111",	-- 0x0FB1
		"11001000",	-- 0x0FB2
		"00001001",	-- 0x0FB3
		"00001001",	-- 0x0FB4
		"01001110",	-- 0x0FB5
		"00100011",	-- 0x0FB6
		"01100110",	-- 0x0FB7
		"01101001",	-- 0x0FB8
		"11101001",	-- 0x0FB9
		"00001010",	-- 0x0FBA
		"00001101",	-- 0x0FBB
		"00001100",	-- 0x0FBC
		"00000111",	-- 0x0FBD
		"00010111",	-- 0x0FBE
		"11001001",	-- 0x0FBF
		"01010101",	-- 0x0FC0
		"11000110",	-- 0x0FC1
		"11111110",	-- 0x0FC2
		"11001000",	-- 0x0FC3
		"00000101",	-- 0x0FC4
		"11001001",	-- 0x0FC5
		"01111001",	-- 0x0FC6
		"11111110",	-- 0x0FC7
		"00100000",	-- 0x0FC8
		"11011010",	-- 0x0FC9
		"10010010",	-- 0x0FCA
		"11000111",	-- 0x0FCB
		"11001011",	-- 0x0FCC
		"10111001",	-- 0x0FCD
		"11001101",	-- 0x0FCE
		"11010100",	-- 0x0FCF
		"11000111",	-- 0x0FD0
		"11000011",	-- 0x0FD1
		"01000010",	-- 0x0FD2
		"11001000",	-- 0x0FD3
		"00101010",	-- 0x0FD4
		"00110110",	-- 0x0FD5
		"11001001",	-- 0x0FD6
		"00000110",	-- 0x0FD7
		"00000000",	-- 0x0FD8
		"00001001",	-- 0x0FD9
		"00001001",	-- 0x0FDA
		"01011110",	-- 0x0FDB
		"00100011",	-- 0x0FDC
		"01100110",	-- 0x0FDD
		"01101011",	-- 0x0FDE
		"00000001",	-- 0x0FDF
		"00001011",	-- 0x0FE0
		"00000000",	-- 0x0FE1
		"00010001",	-- 0x0FE2
		"00001010",	-- 0x0FE3
		"11111100",	-- 0x0FE4
		"11101101",	-- 0x0FE5
		"10110000",	-- 0x0FE6
		"11001101",	-- 0x0FE7
		"11000100",	-- 0x0FE8
		"11000110",	-- 0x0FE9
		"00111110",	-- 0x0FEA
		"01000110",	-- 0x0FEB
		"11010011",	-- 0x0FEC
		"01110001",	-- 0x0FED
		"00111110",	-- 0x0FEE
		"00000001",	-- 0x0FEF
		"00111101",	-- 0x0FF0
		"11010011",	-- 0x0FF1
		"01110000",	-- 0x0FF2
		"00111110",	-- 0x0FF3
		"00110000",	-- 0x0FF4
		"11010011",	-- 0x0FF5
		"01110001",	-- 0x0FF6
		"00011110",	-- 0x0FF7
		"00001001",	-- 0x0FF8
		"00111110",	-- 0x0FF9
		"00010010",	-- 0x0FFA
		"01010111",	-- 0x0FFB
		"11001101",	-- 0x0FFC
		"01111111",	-- 0x0FFD
		"11000111",	-- 0x0FFE
		"00000001");	-- 0x0FFF
begin
	D <= ROM(to_integer(unsigned(A))) when CE_n = '0' and OE_n = '0' else (others => 'Z');
end;
